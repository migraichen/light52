--------------------------------------------------------------------------------
-- obj_code_pkg.vhdl -- Application object code in vhdl constant string format.
--------------------------------------------------------------------------------
-- Written by build_rom.py for project 'Blinker'.
--------------------------------------------------------------------------------
-- Copyright (C) 2012 Jose A. Ruiz
--
-- This source file may be used and distributed without
-- restriction provided that this copyright statement is not
-- removed from the file and that any derivative work contains
-- the original copyright notice and the associated disclaimer.
--
-- This source file is free software; you can redistribute it
-- and/or modify it under the terms of the GNU Lesser General
-- Public License as published by the Free Software Foundation;
-- either version 2.1 of the License, or (at your option) any
-- later version.
--
-- This source is distributed in the hope that it will be
-- useful, but WITHOUT ANY WARRANTY; without even the implied
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
-- PURPOSE.  See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General
-- Public License along with this source; if not, download it
-- from http://www.opencores.org/lgpl.shtml
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.light52_pkg.all;

package obj_code_pkg is

-- Size of XCODE memory in bytes.
constant XCODE_SIZE : natural := 4096;
-- Size of XDATA memory in bytes.
constant XDATA_SIZE : natural := 0;

-- Object code initialization constant.
constant object_code : t_obj_code(0 to 2811) := (
    X"02", X"00", X"11", X"32", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"02", X"01", X"c0", X"02", X"00", 
    X"70", X"75", X"81", X"40", X"12", X"0a", X"b4", X"e5", 
    X"82", X"60", X"03", X"02", X"00", X"0e", X"79", X"00", 
    X"e9", X"44", X"00", X"60", X"1b", X"7a", X"00", X"90", 
    X"0a", X"fc", X"78", X"01", X"75", X"a0", X"00", X"e4", 
    X"93", X"f2", X"a3", X"08", X"b8", X"00", X"02", X"05", 
    X"a0", X"d9", X"f4", X"da", X"f2", X"75", X"a0", X"ff", 
    X"e4", X"78", X"ff", X"f6", X"d8", X"fd", X"78", X"00", 
    X"e8", X"44", X"00", X"60", X"0a", X"79", X"01", X"75", 
    X"a0", X"00", X"e4", X"f3", X"09", X"d8", X"fc", X"78", 
    X"00", X"e8", X"44", X"00", X"60", X"0c", X"79", X"00", 
    X"90", X"00", X"01", X"e4", X"f0", X"a3", X"d8", X"fc", 
    X"d9", X"fa", X"75", X"0c", X"00", X"02", X"00", X"0e", 
    X"12", X"00", X"df", X"74", X"b8", X"c0", X"e0", X"74", 
    X"0a", X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", 
    X"02", X"f6", X"15", X"81", X"15", X"81", X"15", X"81", 
    X"74", X"bb", X"c0", X"e0", X"74", X"0a", X"c0", X"e0", 
    X"74", X"80", X"c0", X"e0", X"12", X"02", X"f6", X"15", 
    X"81", X"15", X"81", X"15", X"81", X"74", X"dd", X"c0", 
    X"e0", X"74", X"0a", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"02", X"f6", X"15", X"81", X"15", X"81", 
    X"15", X"81", X"12", X"01", X"01", X"ac", X"82", X"ad", 
    X"83", X"ae", X"f0", X"ff", X"75", X"37", X"e8", X"75", 
    X"38", X"03", X"e4", X"f5", X"39", X"f5", X"3a", X"8c", 
    X"82", X"8d", X"83", X"8e", X"f0", X"ef", X"12", X"01", 
    X"fb", X"ac", X"82", X"ad", X"83", X"ae", X"f0", X"ff", 
    X"8c", X"90", X"8d", X"80", X"80", X"d4", X"22", X"e4", 
    X"f5", X"08", X"f5", X"09", X"f5", X"0a", X"f5", X"0b", 
    X"90", X"c3", X"50", X"12", X"01", X"6e", X"75", X"82", 
    X"01", X"12", X"01", X"b7", X"75", X"82", X"01", X"12", 
    X"01", X"65", X"75", X"82", X"01", X"12", X"01", X"87", 
    X"22", X"12", X"01", X"90", X"ae", X"82", X"af", X"83", 
    X"7d", X"00", X"7c", X"00", X"75", X"37", X"32", X"e4", 
    X"f5", X"38", X"f5", X"39", X"f5", X"3a", X"8e", X"82", 
    X"8f", X"83", X"8d", X"f0", X"ec", X"12", X"01", X"fb", 
    X"ac", X"82", X"ad", X"83", X"ae", X"f0", X"ff", X"85", 
    X"08", X"37", X"85", X"09", X"38", X"85", X"0a", X"39", 
    X"85", X"0b", X"3a", X"90", X"03", X"e8", X"e4", X"f5", 
    X"f0", X"c0", X"07", X"c0", X"06", X"c0", X"05", X"c0", 
    X"04", X"12", X"02", X"60", X"a8", X"82", X"a9", X"83", 
    X"aa", X"f0", X"fb", X"d0", X"04", X"d0", X"05", X"d0", 
    X"06", X"d0", X"07", X"e8", X"2c", X"fc", X"e9", X"3d", 
    X"fd", X"ea", X"3e", X"fe", X"eb", X"3f", X"8c", X"82", 
    X"8d", X"83", X"8e", X"f0", X"22", X"e5", X"82", X"54", 
    X"01", X"24", X"ff", X"92", X"af", X"22", X"ae", X"82", 
    X"af", X"83", X"be", X"ff", X"05", X"bf", X"ff", X"02", 
    X"80", X"08", X"8f", X"8f", X"8e", X"8e", X"d2", X"8c", 
    X"80", X"02", X"c2", X"8c", X"d2", X"88", X"22", X"e5", 
    X"82", X"54", X"01", X"24", X"ff", X"92", X"8d", X"22", 
    X"85", X"8d", X"37", X"85", X"8c", X"38", X"85", X"8c", 
    X"39", X"e5", X"39", X"b5", X"38", X"02", X"80", X"06", 
    X"85", X"8d", X"37", X"85", X"8c", X"38", X"af", X"37", 
    X"7e", X"00", X"ac", X"38", X"7d", X"00", X"ec", X"4e", 
    X"f5", X"82", X"ed", X"4f", X"f5", X"83", X"22", X"e5", 
    X"82", X"54", X"01", X"24", X"ff", X"92", X"a9", X"22", 
    X"c0", X"e0", X"c0", X"d0", X"d2", X"88", X"85", X"0c", 
    X"90", X"05", X"0c", X"74", X"01", X"25", X"08", X"f5", 
    X"08", X"e4", X"35", X"09", X"f5", X"09", X"e4", X"35", 
    X"0a", X"f5", X"0a", X"e4", X"35", X"0b", X"f5", X"0b", 
    X"d0", X"d0", X"d0", X"e0", X"32", X"ae", X"82", X"af", 
    X"83", X"30", X"9c", X"fd", X"8e", X"99", X"be", X"0a", 
    X"09", X"bf", X"00", X"06", X"30", X"9c", X"fd", X"75", 
    X"99", X"0d", X"22", X"fb", X"7a", X"20", X"e4", X"fc", 
    X"fd", X"fe", X"ff", X"e5", X"82", X"25", X"82", X"f5", 
    X"82", X"e5", X"83", X"33", X"f5", X"83", X"e5", X"f0", 
    X"33", X"f5", X"f0", X"eb", X"33", X"fb", X"40", X"17", 
    X"da", X"e9", X"80", X"42", X"e5", X"82", X"25", X"82", 
    X"f5", X"82", X"e5", X"83", X"33", X"f5", X"83", X"e5", 
    X"f0", X"33", X"f5", X"f0", X"eb", X"33", X"fb", X"ec", 
    X"33", X"fc", X"ed", X"33", X"fd", X"ee", X"33", X"fe", 
    X"ef", X"33", X"ff", X"ec", X"95", X"37", X"ed", X"95", 
    X"38", X"ee", X"95", X"39", X"ef", X"95", X"3a", X"40", 
    X"13", X"ec", X"95", X"37", X"fc", X"ed", X"95", X"38", 
    X"fd", X"ee", X"95", X"39", X"fe", X"ef", X"95", X"3a", 
    X"ff", X"43", X"82", X"01", X"da", X"be", X"eb", X"22", 
    X"aa", X"f0", X"fb", X"e5", X"82", X"85", X"37", X"f0", 
    X"a4", X"fc", X"ad", X"f0", X"e5", X"83", X"85", X"37", 
    X"f0", X"a4", X"2d", X"fd", X"e4", X"35", X"f0", X"fe", 
    X"e5", X"82", X"85", X"38", X"f0", X"a4", X"2d", X"fd", 
    X"e5", X"f0", X"3e", X"fe", X"e4", X"33", X"ff", X"ea", 
    X"85", X"37", X"f0", X"a4", X"2e", X"fe", X"e5", X"f0", 
    X"3f", X"ff", X"e5", X"83", X"85", X"38", X"f0", X"a4", 
    X"2e", X"fe", X"e5", X"f0", X"3f", X"ff", X"e5", X"82", 
    X"85", X"39", X"f0", X"a4", X"2e", X"fe", X"e5", X"f0", 
    X"3f", X"ff", X"eb", X"85", X"37", X"f0", X"a4", X"2f", 
    X"ff", X"ea", X"85", X"38", X"f0", X"a4", X"2f", X"ff", 
    X"e5", X"83", X"85", X"39", X"f0", X"a4", X"2f", X"ff", 
    X"e5", X"82", X"85", X"3a", X"f0", X"a4", X"2f", X"8e", 
    X"f0", X"8d", X"83", X"8c", X"82", X"22", X"c0", X"36", 
    X"85", X"81", X"36", X"7e", X"00", X"8e", X"83", X"12", 
    X"01", X"e5", X"d0", X"36", X"22", X"85", X"82", X"1e", 
    X"85", X"83", X"1f", X"85", X"f0", X"20", X"e4", X"f5", 
    X"1b", X"f5", X"1c", X"f5", X"1d", X"85", X"0d", X"21", 
    X"90", X"02", X"ce", X"02", X"03", X"c3", X"c0", X"36", 
    X"85", X"81", X"36", X"e5", X"36", X"24", X"fb", X"ff", 
    X"8f", X"21", X"e4", X"f5", X"1b", X"f5", X"1c", X"f5", 
    X"1d", X"e5", X"36", X"24", X"fb", X"f8", X"86", X"1e", 
    X"08", X"86", X"1f", X"08", X"86", X"20", X"90", X"02", 
    X"ce", X"12", X"03", X"c3", X"d0", X"36", X"22", X"af", 
    X"82", X"c0", X"11", X"c0", X"12", X"c0", X"13", X"12", 
    X"03", X"2c", X"80", X"07", X"c0", X"0f", X"c0", X"10", 
    X"8f", X"82", X"22", X"15", X"81", X"15", X"81", X"15", 
    X"81", X"05", X"19", X"e4", X"b5", X"19", X"02", X"05", 
    X"1a", X"22", X"af", X"82", X"74", X"30", X"2f", X"ff", 
    X"24", X"c6", X"50", X"11", X"74", X"07", X"2f", X"ff", 
    X"e5", X"0e", X"60", X"09", X"8f", X"05", X"7e", X"00", 
    X"43", X"05", X"20", X"8d", X"07", X"8f", X"82", X"02", 
    X"03", X"1f", X"e5", X"82", X"ff", X"c4", X"54", X"0f", 
    X"f5", X"82", X"c0", X"07", X"12", X"03", X"42", X"d0", 
    X"07", X"74", X"0f", X"5f", X"f5", X"82", X"02", X"03", 
    X"42", X"85", X"82", X"37", X"ab", X"14", X"ac", X"15", 
    X"ad", X"16", X"ae", X"17", X"aa", X"18", X"75", X"39", 
    X"20", X"8a", X"07", X"ef", X"2f", X"f5", X"38", X"ee", 
    X"23", X"54", X"01", X"45", X"38", X"fa", X"eb", X"2b", 
    X"fb", X"ec", X"33", X"fc", X"ed", X"33", X"fd", X"ee", 
    X"33", X"fe", X"c3", X"ea", X"95", X"37", X"40", X"08", 
    X"ea", X"c3", X"95", X"37", X"fa", X"43", X"03", X"01", 
    X"e5", X"39", X"14", X"ff", X"8f", X"39", X"70", X"d1", 
    X"8b", X"14", X"8c", X"15", X"8d", X"16", X"8e", X"17", 
    X"8a", X"18", X"22", X"85", X"82", X"0f", X"85", X"83", 
    X"10", X"85", X"1b", X"11", X"85", X"1c", X"12", X"85", 
    X"1d", X"13", X"e4", X"f5", X"19", X"f5", X"1a", X"ad", 
    X"1e", X"ae", X"1f", X"af", X"20", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"0a", X"98", X"fc", X"74", 
    X"01", X"2d", X"f5", X"1e", X"e4", X"3e", X"f5", X"1f", 
    X"8f", X"20", X"ec", X"ff", X"70", X"03", X"02", X"0a", 
    X"79", X"bf", X"25", X"02", X"80", X"03", X"02", X"0a", 
    X"71", X"7e", X"00", X"7d", X"00", X"8e", X"22", X"8e", 
    X"23", X"7a", X"00", X"7b", X"00", X"8e", X"24", X"7c", 
    X"00", X"8e", X"25", X"8e", X"2b", X"75", X"26", X"ff", 
    X"85", X"1e", X"2c", X"85", X"1f", X"2d", X"85", X"20", 
    X"2e", X"85", X"2c", X"82", X"85", X"2d", X"83", X"85", 
    X"2e", X"f0", X"12", X"0a", X"98", X"f5", X"2f", X"a3", 
    X"85", X"82", X"2c", X"85", X"83", X"2d", X"85", X"2c", 
    X"1e", X"85", X"2d", X"1f", X"85", X"2e", X"20", X"74", 
    X"25", X"b5", X"2f", X"08", X"85", X"2f", X"82", X"12", 
    X"03", X"1f", X"80", X"8b", X"74", X"d0", X"25", X"2f", 
    X"50", X"39", X"e5", X"2f", X"24", X"c6", X"40", X"33", 
    X"74", X"ff", X"b5", X"26", X"1a", X"e5", X"2b", X"f5", 
    X"30", X"75", X"f0", X"0a", X"a4", X"f5", X"30", X"e5", 
    X"2f", X"f5", X"31", X"25", X"30", X"24", X"d0", X"f5", 
    X"2b", X"70", X"ae", X"7d", X"01", X"80", X"aa", X"e5", 
    X"26", X"75", X"f0", X"0a", X"a4", X"f5", X"31", X"e5", 
    X"2f", X"f5", X"30", X"25", X"31", X"24", X"d0", X"f5", 
    X"26", X"80", X"96", X"74", X"2e", X"b5", X"2f", X"0a", 
    X"74", X"ff", X"b5", X"26", X"8c", X"75", X"26", X"00", 
    X"80", X"87", X"74", X"9f", X"25", X"2f", X"50", X"0e", 
    X"e5", X"2f", X"24", X"85", X"40", X"08", X"53", X"2f", 
    X"df", X"75", X"0e", X"01", X"80", X"03", X"75", X"0e", 
    X"00", X"74", X"20", X"b5", X"2f", X"03", X"02", X"05", 
    X"4c", X"74", X"2b", X"b5", X"2f", X"03", X"02", X"05", 
    X"46", X"74", X"2d", X"b5", X"2f", X"02", X"80", X"79", 
    X"74", X"42", X"b5", X"2f", X"03", X"02", X"05", X"52", 
    X"74", X"43", X"b5", X"2f", X"03", X"02", X"05", X"5d", 
    X"74", X"44", X"b5", X"2f", X"03", X"02", X"07", X"6e", 
    X"74", X"46", X"b5", X"2f", X"03", X"02", X"07", X"84", 
    X"74", X"48", X"b5", X"2f", X"03", X"02", X"04", X"21", 
    X"74", X"49", X"b5", X"2f", X"03", X"02", X"07", X"6e", 
    X"74", X"4a", X"b5", X"2f", X"03", X"02", X"04", X"21", 
    X"74", X"4c", X"b5", X"2f", X"02", X"80", X"50", X"74", 
    X"4f", X"b5", X"2f", X"03", X"02", X"07", X"75", X"74", 
    X"50", X"b5", X"2f", X"03", X"02", X"06", X"b9", X"74", 
    X"53", X"b5", X"2f", X"02", X"80", X"76", X"74", X"54", 
    X"b5", X"2f", X"03", X"02", X"04", X"21", X"74", X"55", 
    X"b5", X"2f", X"03", X"02", X"07", X"7a", X"74", X"58", 
    X"b5", X"2f", X"03", X"02", X"07", X"7f", X"74", X"5a", 
    X"b5", X"2f", X"03", X"02", X"04", X"21", X"02", X"07", 
    X"88", X"7e", X"01", X"02", X"04", X"21", X"75", X"22", 
    X"01", X"02", X"04", X"21", X"75", X"23", X"01", X"02", 
    X"04", X"21", X"7b", X"01", X"02", X"04", X"21", X"75", 
    X"24", X"01", X"02", X"04", X"21", X"eb", X"60", X"0a", 
    X"e5", X"21", X"14", X"f9", X"89", X"21", X"87", X"31", 
    X"80", X"0d", X"e5", X"21", X"24", X"fe", X"f5", X"30", 
    X"85", X"30", X"21", X"a9", X"30", X"87", X"31", X"85", 
    X"31", X"82", X"c0", X"06", X"c0", X"05", X"c0", X"04", 
    X"c0", X"03", X"c0", X"02", X"12", X"03", X"1f", X"d0", 
    X"02", X"d0", X"03", X"d0", X"04", X"d0", X"05", X"d0", 
    X"06", X"02", X"07", X"a7", X"e5", X"21", X"24", X"fd", 
    X"f5", X"31", X"85", X"31", X"21", X"a9", X"31", X"87", 
    X"2c", X"09", X"87", X"2d", X"09", X"87", X"2e", X"19", 
    X"19", X"85", X"2c", X"14", X"85", X"2d", X"15", X"85", 
    X"2e", X"16", X"85", X"2c", X"82", X"85", X"2d", X"83", 
    X"85", X"2e", X"f0", X"c0", X"06", X"c0", X"05", X"c0", 
    X"04", X"c0", X"03", X"c0", X"02", X"12", X"0a", X"80", 
    X"85", X"82", X"2c", X"85", X"83", X"2d", X"d0", X"02", 
    X"d0", X"03", X"d0", X"04", X"d0", X"05", X"d0", X"06", 
    X"85", X"2c", X"31", X"74", X"ff", X"b5", X"26", X"03", 
    X"85", X"31", X"26", X"ee", X"70", X"36", X"c3", X"e5", 
    X"31", X"95", X"2b", X"50", X"2f", X"e5", X"2b", X"c3", 
    X"95", X"31", X"f5", X"30", X"85", X"30", X"2c", X"15", 
    X"30", X"e5", X"2c", X"60", X"1c", X"75", X"82", X"20", 
    X"c0", X"06", X"c0", X"05", X"c0", X"04", X"c0", X"03", 
    X"c0", X"02", X"12", X"03", X"1f", X"d0", X"02", X"d0", 
    X"03", X"d0", X"04", X"d0", X"05", X"d0", X"06", X"80", 
    X"db", X"85", X"30", X"2b", X"85", X"26", X"30", X"85", 
    X"14", X"82", X"85", X"15", X"83", X"85", X"16", X"f0", 
    X"12", X"0a", X"98", X"f5", X"2c", X"85", X"2c", X"28", 
    X"60", X"48", X"85", X"30", X"2c", X"15", X"30", X"c3", 
    X"74", X"80", X"85", X"2c", X"f0", X"63", X"f0", X"80", 
    X"95", X"f0", X"50", X"36", X"85", X"28", X"82", X"c0", 
    X"06", X"c0", X"05", X"c0", X"04", X"c0", X"03", X"c0", 
    X"02", X"12", X"03", X"1f", X"d0", X"02", X"d0", X"03", 
    X"d0", X"04", X"d0", X"05", X"d0", X"06", X"85", X"14", 
    X"2c", X"85", X"15", X"2d", X"85", X"16", X"2e", X"05", 
    X"2c", X"e4", X"b5", X"2c", X"02", X"05", X"2d", X"85", 
    X"2c", X"14", X"85", X"2d", X"15", X"85", X"2e", X"16", 
    X"80", X"a5", X"ee", X"70", X"03", X"02", X"07", X"a7", 
    X"c3", X"e5", X"31", X"95", X"2b", X"40", X"03", X"02", 
    X"07", X"a7", X"e5", X"2b", X"c3", X"95", X"31", X"f5", 
    X"31", X"85", X"31", X"30", X"15", X"31", X"e5", X"30", 
    X"70", X"03", X"02", X"07", X"a4", X"75", X"82", X"20", 
    X"c0", X"06", X"c0", X"05", X"c0", X"04", X"c0", X"03", 
    X"c0", X"02", X"12", X"03", X"1f", X"d0", X"02", X"d0", 
    X"03", X"d0", X"04", X"d0", X"05", X"d0", X"06", X"80", 
    X"d8", X"e5", X"21", X"24", X"fd", X"f5", X"30", X"85", 
    X"30", X"21", X"a9", X"30", X"87", X"2c", X"09", X"87", 
    X"2d", X"09", X"87", X"2e", X"19", X"19", X"85", X"2c", 
    X"14", X"85", X"2d", X"15", X"85", X"2e", X"16", X"85", 
    X"16", X"29", X"74", X"80", X"25", X"29", X"50", X"05", 
    X"75", X"30", X"43", X"80", X"19", X"74", X"a0", X"25", 
    X"29", X"50", X"05", X"75", X"30", X"50", X"80", X"0e", 
    X"74", X"c0", X"25", X"29", X"50", X"05", X"75", X"30", 
    X"49", X"80", X"03", X"75", X"30", X"58", X"85", X"30", 
    X"82", X"c0", X"06", X"c0", X"05", X"c0", X"04", X"c0", 
    X"03", X"c0", X"02", X"12", X"03", X"1f", X"75", X"82", 
    X"3a", X"12", X"03", X"1f", X"75", X"82", X"30", X"12", 
    X"03", X"1f", X"75", X"82", X"78", X"12", X"03", X"1f", 
    X"d0", X"02", X"d0", X"03", X"d0", X"04", X"d0", X"05", 
    X"d0", X"06", X"74", X"49", X"b5", X"30", X"02", X"80", 
    X"21", X"74", X"50", X"b5", X"30", X"02", X"80", X"1a", 
    X"85", X"15", X"82", X"c0", X"06", X"c0", X"05", X"c0", 
    X"04", X"c0", X"03", X"c0", X"02", X"12", X"03", X"62", 
    X"d0", X"02", X"d0", X"03", X"d0", X"04", X"d0", X"05", 
    X"d0", X"06", X"85", X"14", X"82", X"c0", X"06", X"c0", 
    X"05", X"c0", X"04", X"c0", X"03", X"c0", X"02", X"12", 
    X"03", X"62", X"d0", X"02", X"d0", X"03", X"d0", X"04", 
    X"d0", X"05", X"d0", X"06", X"80", X"39", X"7a", X"01", 
    X"75", X"25", X"0a", X"80", X"32", X"75", X"25", X"08", 
    X"80", X"2d", X"75", X"25", X"0a", X"80", X"28", X"75", 
    X"25", X"10", X"80", X"23", X"7c", X"01", X"80", X"1f", 
    X"85", X"2f", X"82", X"c0", X"06", X"c0", X"05", X"c0", 
    X"04", X"c0", X"03", X"c0", X"02", X"12", X"03", X"1f", 
    X"d0", X"02", X"d0", X"03", X"d0", X"04", X"d0", X"05", 
    X"d0", X"06", X"80", X"03", X"85", X"31", X"2b", X"ec", 
    X"60", X"68", X"e5", X"21", X"24", X"fc", X"fc", X"8c", 
    X"21", X"8c", X"01", X"87", X"32", X"09", X"87", X"33", 
    X"09", X"87", X"34", X"09", X"87", X"35", X"19", X"19", 
    X"19", X"85", X"32", X"14", X"85", X"33", X"15", X"85", 
    X"34", X"16", X"85", X"35", X"17", X"75", X"14", X"f1", 
    X"75", X"15", X"0a", X"75", X"16", X"80", X"85", X"14", 
    X"32", X"85", X"15", X"33", X"85", X"16", X"34", X"74", 
    X"01", X"25", X"32", X"f5", X"2c", X"e4", X"35", X"33", 
    X"f5", X"2d", X"85", X"34", X"2e", X"85", X"2c", X"14", 
    X"85", X"2d", X"15", X"85", X"2e", X"16", X"85", X"32", 
    X"82", X"85", X"33", X"83", X"85", X"34", X"f0", X"12", 
    X"0a", X"98", X"fc", X"8c", X"32", X"70", X"03", X"02", 
    X"03", X"d7", X"85", X"32", X"82", X"12", X"03", X"1f", 
    X"80", X"c4", X"e5", X"25", X"70", X"03", X"02", X"03", 
    X"d7", X"eb", X"60", X"3f", X"e5", X"21", X"14", X"f9", 
    X"89", X"21", X"87", X"04", X"8c", X"32", X"75", X"33", 
    X"00", X"75", X"34", X"00", X"75", X"35", X"00", X"85", 
    X"32", X"14", X"85", X"33", X"15", X"85", X"34", X"16", 
    X"85", X"35", X"17", X"ea", X"60", X"03", X"02", X"08", 
    X"c4", X"85", X"14", X"32", X"75", X"33", X"00", X"75", 
    X"34", X"00", X"75", X"35", X"00", X"85", X"32", X"14", 
    X"85", X"33", X"15", X"85", X"34", X"16", X"85", X"35", 
    X"17", X"80", X"69", X"e5", X"24", X"60", X"25", X"e5", 
    X"21", X"24", X"fc", X"fc", X"8c", X"21", X"8c", X"01", 
    X"87", X"32", X"09", X"87", X"33", X"09", X"87", X"34", 
    X"09", X"87", X"35", X"19", X"19", X"19", X"85", X"32", 
    X"14", X"85", X"33", X"15", X"85", X"34", X"16", X"85", 
    X"35", X"17", X"80", X"40", X"e5", X"21", X"24", X"fe", 
    X"fc", X"8c", X"21", X"8c", X"01", X"87", X"03", X"09", 
    X"87", X"04", X"19", X"8b", X"32", X"ec", X"f5", X"33", 
    X"33", X"95", X"e0", X"f5", X"34", X"f5", X"35", X"85", 
    X"32", X"14", X"85", X"33", X"15", X"85", X"34", X"16", 
    X"85", X"35", X"17", X"ea", X"70", X"16", X"85", X"14", 
    X"32", X"85", X"15", X"33", X"f5", X"34", X"f5", X"35", 
    X"85", X"32", X"14", X"85", X"33", X"15", X"85", X"34", 
    X"16", X"85", X"35", X"17", X"ea", X"60", X"2a", X"e5", 
    X"17", X"30", X"e7", X"23", X"c3", X"e4", X"95", X"14", 
    X"f5", X"32", X"e4", X"95", X"15", X"f5", X"33", X"e4", 
    X"95", X"16", X"f5", X"34", X"e4", X"95", X"17", X"f5", 
    X"35", X"85", X"32", X"14", X"85", X"33", X"15", X"85", 
    X"34", X"16", X"85", X"35", X"17", X"80", X"02", X"7a", 
    X"00", X"7c", X"01", X"79", X"40", X"7b", X"00", X"75", 
    X"18", X"00", X"85", X"25", X"82", X"c0", X"06", X"c0", 
    X"05", X"c0", X"04", X"c0", X"03", X"c0", X"02", X"c0", 
    X"01", X"12", X"03", X"79", X"d0", X"01", X"d0", X"02", 
    X"d0", X"03", X"d0", X"04", X"d0", X"05", X"d0", X"06", 
    X"ec", X"70", X"10", X"c0", X"03", X"e5", X"18", X"c4", 
    X"f5", X"32", X"e7", X"45", X"32", X"f7", X"19", X"d0", 
    X"03", X"80", X"02", X"a7", X"18", X"0b", X"ec", X"b4", 
    X"01", X"00", X"e4", X"33", X"fc", X"e5", X"14", X"45", 
    X"15", X"45", X"16", X"45", X"17", X"70", X"b8", X"89", 
    X"2a", X"8b", X"27", X"e5", X"2b", X"70", X"03", X"75", 
    X"2b", X"01", X"ed", X"70", X"2c", X"ee", X"70", X"29", 
    X"85", X"2b", X"32", X"ab", X"27", X"0b", X"c3", X"eb", 
    X"95", X"32", X"50", X"1a", X"75", X"82", X"20", X"c0", 
    X"06", X"c0", X"05", X"c0", X"04", X"c0", X"02", X"12", 
    X"03", X"1f", X"d0", X"02", X"d0", X"04", X"d0", X"05", 
    X"d0", X"06", X"15", X"32", X"80", X"dd", X"85", X"32", 
    X"2b", X"ea", X"60", X"16", X"75", X"82", X"2d", X"c0", 
    X"06", X"c0", X"05", X"c0", X"04", X"12", X"03", X"1f", 
    X"d0", X"04", X"d0", X"05", X"d0", X"06", X"15", X"2b", 
    X"80", X"36", X"e5", X"27", X"60", X"32", X"e5", X"22", 
    X"60", X"16", X"75", X"82", X"2b", X"c0", X"06", X"c0", 
    X"05", X"c0", X"04", X"12", X"03", X"1f", X"d0", X"04", 
    X"d0", X"05", X"d0", X"06", X"15", X"2b", X"80", X"18", 
    X"e5", X"23", X"60", X"14", X"75", X"82", X"20", X"c0", 
    X"06", X"c0", X"05", X"c0", X"04", X"12", X"03", X"1f", 
    X"d0", X"04", X"d0", X"05", X"d0", X"06", X"15", X"2b", 
    X"ee", X"70", X"34", X"ab", X"2b", X"8b", X"02", X"1b", 
    X"c3", X"e5", X"27", X"9a", X"50", X"3c", X"ed", X"60", 
    X"08", X"75", X"32", X"30", X"75", X"33", X"00", X"80", 
    X"06", X"75", X"32", X"20", X"75", X"33", X"00", X"85", 
    X"32", X"82", X"c0", X"06", X"c0", X"05", X"c0", X"04", 
    X"c0", X"03", X"12", X"03", X"1f", X"d0", X"03", X"d0", 
    X"04", X"d0", X"05", X"d0", X"06", X"80", X"ce", X"c3", 
    X"e5", X"27", X"95", X"2b", X"50", X"08", X"e5", X"2b", 
    X"c3", X"95", X"27", X"fd", X"80", X"06", X"7d", X"00", 
    X"80", X"02", X"8b", X"05", X"a9", X"2a", X"ab", X"27", 
    X"8b", X"02", X"1b", X"ea", X"60", X"36", X"ec", X"b4", 
    X"01", X"00", X"e4", X"33", X"fc", X"70", X"0a", X"09", 
    X"e7", X"c4", X"54", X"0f", X"fa", X"8a", X"18", X"80", 
    X"07", X"87", X"02", X"74", X"0f", X"5a", X"f5", X"18", 
    X"85", X"18", X"82", X"c0", X"06", X"c0", X"05", X"c0", 
    X"04", X"c0", X"03", X"c0", X"01", X"12", X"03", X"42", 
    X"d0", X"01", X"d0", X"03", X"d0", X"04", X"d0", X"05", 
    X"d0", X"06", X"80", X"c4", X"ee", X"70", X"03", X"02", 
    X"03", X"d7", X"8d", X"06", X"8e", X"05", X"1e", X"ed", 
    X"70", X"03", X"02", X"03", X"d7", X"75", X"82", X"20", 
    X"c0", X"06", X"12", X"03", X"1f", X"d0", X"06", X"80", 
    X"eb", X"8f", X"82", X"12", X"03", X"1f", X"02", X"03", 
    X"d7", X"85", X"19", X"82", X"85", X"1a", X"83", X"22", 
    X"aa", X"82", X"ab", X"83", X"12", X"0a", X"98", X"60", 
    X"03", X"a3", X"80", X"f8", X"c3", X"e5", X"82", X"9a", 
    X"f5", X"82", X"e5", X"83", X"9b", X"f5", X"83", X"22", 
    X"20", X"f7", X"14", X"30", X"f6", X"14", X"88", X"83", 
    X"a8", X"82", X"20", X"f5", X"07", X"e6", X"a8", X"83", 
    X"75", X"83", X"00", X"22", X"e2", X"80", X"f7", X"e4", 
    X"93", X"22", X"e0", X"22", X"75", X"82", X"00", X"22", 
    X"0a", X"0d", X"00", X"4c", X"69", X"67", X"68", X"74", 
    X"35", X"32", X"20", X"70", X"72", X"6f", X"6a", X"65", 
    X"63", X"74", X"20", X"2d", X"2d", X"20", X"41", X"75", 
    X"67", X"20", X"32", X"30", X"20", X"32", X"30", X"31", 
    X"38", X"0a", X"0a", X"0d", X"00", X"4c", X"45", X"44", 
    X"20", X"62", X"6c", X"69", X"6e", X"6b", X"65", X"72", 
    X"20", X"74", X"65", X"73", X"74", X"2e", X"0a", X"0d", 
    X"00", X"3c", X"4e", X"4f", X"20", X"46", X"4c", X"4f", 
    X"41", X"54", X"3e", X"00" 
);


end package obj_code_pkg;

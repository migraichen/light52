--------------------------------------------------------------------------------
-- obj_code_pkg.vhdl -- Application object code in vhdl constant string format.
--------------------------------------------------------------------------------
-- Written by build_rom.py for project 'FreeRTOS'.
--------------------------------------------------------------------------------
-- Copyright (C) 2012 Jose A. Ruiz
--
-- This source file may be used and distributed without
-- restriction provided that this copyright statement is not
-- removed from the file and that any derivative work contains
-- the original copyright notice and the associated disclaimer.
--
-- This source file is free software; you can redistribute it
-- and/or modify it under the terms of the GNU Lesser General
-- Public License as published by the Free Software Foundation;
-- either version 2.1 of the License, or (at your option) any
-- later version.
--
-- This source is distributed in the hope that it will be
-- useful, but WITHOUT ANY WARRANTY; without even the implied
-- warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR
-- PURPOSE.  See the GNU Lesser General Public License for more
-- details.
--
-- You should have received a copy of the GNU Lesser General
-- Public License along with this source; if not, download it
-- from http://www.opencores.org/lgpl.shtml
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.light52_pkg.all;

package obj_code_pkg is

-- Size of XCODE memory in bytes.
constant XCODE_SIZE : natural := 32768;
-- Size of XDATA memory in bytes.
constant XDATA_SIZE : natural := 8192;

-- Object code initialization constant.
constant object_code : t_obj_code(0 to 28922) := (
    X"02", X"00", X"3f", X"32", X"00", X"00", X"00", X"00", 
    X"00", X"00", X"00", X"02", X"65", X"91", X"02", X"00", 
    X"c5", X"e5", X"81", X"24", X"fc", X"c3", X"c8", X"c0", 
    X"e0", X"c0", X"82", X"e6", X"08", X"46", X"70", X"06", 
    X"e5", X"82", X"45", X"83", X"60", X"12", X"18", X"e5", 
    X"82", X"96", X"f5", X"82", X"08", X"e5", X"83", X"96", 
    X"42", X"82", X"08", X"e5", X"f0", X"96", X"45", X"82", 
    X"d0", X"82", X"c8", X"d0", X"e0", X"c8", X"22", X"75", 
    X"81", X"20", X"12", X"70", X"76", X"e5", X"82", X"60", 
    X"03", X"02", X"00", X"0e", X"e4", X"78", X"7f", X"f6", 
    X"d8", X"fd", X"90", X"00", X"03", X"74", X"7a", X"f0", 
    X"74", X"70", X"a3", X"f0", X"74", X"80", X"a3", X"f0", 
    X"90", X"00", X"06", X"74", X"81", X"f0", X"74", X"70", 
    X"a3", X"f0", X"74", X"80", X"a3", X"f0", X"90", X"00", 
    X"01", X"e4", X"f0", X"a3", X"f0", X"90", X"00", X"09", 
    X"e4", X"f0", X"a3", X"f0", X"a3", X"f0", X"90", X"00", 
    X"66", X"f0", X"90", X"00", X"67", X"f0", X"a3", X"f0", 
    X"90", X"00", X"69", X"f0", X"90", X"00", X"6a", X"f0", 
    X"90", X"00", X"6b", X"f0", X"90", X"00", X"6c", X"f0", 
    X"90", X"00", X"6d", X"f0", X"90", X"00", X"6e", X"f0", 
    X"90", X"00", X"6f", X"f0", X"a3", X"f0", X"90", X"00", 
    X"71", X"f0", X"a3", X"f0", X"a3", X"f0", X"90", X"00", 
    X"74", X"f0", X"90", X"18", X"77", X"e4", X"f0", X"a3", 
    X"f0", X"a3", X"f0", X"90", X"18", X"75", X"e4", X"f0", 
    X"a3", X"f0", X"02", X"00", X"0e", X"12", X"01", X"83", 
    X"74", X"88", X"c0", X"e0", X"74", X"70", X"c0", X"e0", 
    X"74", X"80", X"c0", X"e0", X"12", X"67", X"c5", X"15", 
    X"81", X"15", X"81", X"15", X"81", X"74", X"8b", X"c0", 
    X"e0", X"74", X"70", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"12", X"67", X"c5", X"15", X"81", X"15", X"81", 
    X"15", X"81", X"74", X"b6", X"c0", X"e0", X"74", X"70", 
    X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", X"67", 
    X"c5", X"15", X"81", X"15", X"81", X"15", X"81", X"90", 
    X"00", X"03", X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", 
    X"e0", X"ff", X"e4", X"c0", X"e0", X"c0", X"e0", X"c0", 
    X"e0", X"04", X"c0", X"e0", X"c0", X"05", X"c0", X"06", 
    X"c0", X"07", X"74", X"e8", X"c0", X"e0", X"74", X"03", 
    X"c0", X"e0", X"74", X"c7", X"c0", X"e0", X"74", X"70", 
    X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"90", X"01", 
    X"8a", X"12", X"02", X"80", X"e5", X"81", X"24", X"f4", 
    X"f5", X"81", X"90", X"00", X"06", X"e0", X"fd", X"a3", 
    X"e0", X"fe", X"a3", X"e0", X"ff", X"e4", X"c0", X"e0", 
    X"c0", X"e0", X"c0", X"e0", X"04", X"c0", X"e0", X"c0", 
    X"05", X"c0", X"06", X"c0", X"07", X"74", X"e8", X"c0", 
    X"e0", X"74", X"03", X"c0", X"e0", X"74", X"d1", X"c0", 
    X"e0", X"74", X"70", X"c0", X"e0", X"74", X"80", X"c0", 
    X"e0", X"90", X"02", X"16", X"12", X"02", X"80", X"e5", 
    X"81", X"24", X"f4", X"f5", X"81", X"12", X"08", X"ed", 
    X"80", X"fe", X"22", X"75", X"80", X"00", X"75", X"90", 
    X"00", X"22", X"ad", X"82", X"ae", X"83", X"af", X"f0", 
    X"90", X"00", X"01", X"e0", X"f5", X"f0", X"a3", X"e0", 
    X"45", X"f0", X"70", X"f4", X"90", X"00", X"01", X"74", 
    X"01", X"f0", X"e4", X"a3", X"f0", X"c0", X"05", X"c0", 
    X"06", X"c0", X"07", X"74", X"d8", X"c0", X"e0", X"74", 
    X"70", X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", 
    X"67", X"c5", X"e5", X"81", X"24", X"fa", X"f5", X"81", 
    X"90", X"00", X"01", X"e4", X"f0", X"a3", X"f0", X"90", 
    X"00", X"01", X"e0", X"f5", X"f0", X"a3", X"e0", X"45", 
    X"f0", X"70", X"f4", X"90", X"00", X"01", X"74", X"01", 
    X"f0", X"e4", X"a3", X"f0", X"74", X"57", X"c0", X"e0", 
    X"e4", X"c0", X"e0", X"74", X"e8", X"c0", X"e0", X"74", 
    X"70", X"c0", X"e0", X"74", X"80", X"c0", X"e0", X"12", 
    X"67", X"c5", X"e5", X"81", X"24", X"fb", X"f5", X"81", 
    X"90", X"00", X"01", X"e4", X"f0", X"a3", X"f0", X"ae", 
    X"80", X"63", X"06", X"ff", X"8e", X"80", X"ae", X"90", 
    X"63", X"06", X"ff", X"8e", X"90", X"90", X"00", X"64", 
    X"12", X"08", X"be", X"80", X"b2", X"22", X"ad", X"82", 
    X"ae", X"83", X"af", X"f0", X"90", X"00", X"01", X"e0", 
    X"f5", X"f0", X"a3", X"e0", X"45", X"f0", X"70", X"f4", 
    X"90", X"00", X"01", X"74", X"01", X"f0", X"e4", X"a3", 
    X"f0", X"c0", X"05", X"c0", X"06", X"c0", X"07", X"74", 
    X"d8", X"c0", X"e0", X"74", X"70", X"c0", X"e0", X"74", 
    X"80", X"c0", X"e0", X"12", X"67", X"c5", X"e5", X"81", 
    X"24", X"fa", X"f5", X"81", X"90", X"00", X"01", X"e4", 
    X"f0", X"a3", X"f0", X"12", X"66", X"98", X"ae", X"82", 
    X"90", X"00", X"01", X"e0", X"f5", X"f0", X"a3", X"e0", 
    X"45", X"f0", X"70", X"f4", X"90", X"00", X"01", X"74", 
    X"01", X"f0", X"e4", X"a3", X"f0", X"7f", X"00", X"8e", 
    X"82", X"8f", X"83", X"12", X"66", X"87", X"90", X"00", 
    X"01", X"e4", X"f0", X"a3", X"f0", X"80", X"d4", X"22", 
    X"c0", X"0c", X"85", X"81", X"0c", X"05", X"81", X"05", 
    X"81", X"05", X"81", X"ae", X"82", X"af", X"83", X"90", 
    X"00", X"33", X"c0", X"07", X"c0", X"06", X"12", X"61", 
    X"84", X"ab", X"82", X"ac", X"83", X"ad", X"f0", X"d0", 
    X"06", X"d0", X"07", X"a8", X"0c", X"08", X"a6", X"03", 
    X"08", X"a6", X"04", X"08", X"a6", X"05", X"a8", X"0c", 
    X"08", X"e6", X"08", X"46", X"60", X"77", X"c0", X"06", 
    X"c0", X"07", X"a8", X"0c", X"08", X"74", X"20", X"26", 
    X"fa", X"e4", X"08", X"36", X"fe", X"08", X"86", X"07", 
    X"e5", X"0c", X"24", X"f9", X"f8", X"86", X"04", X"08", 
    X"86", X"05", X"8c", X"82", X"8d", X"83", X"c0", X"07", 
    X"c0", X"06", X"c0", X"02", X"12", X"61", X"84", X"ab", 
    X"82", X"ac", X"83", X"ad", X"f0", X"d0", X"02", X"d0", 
    X"06", X"d0", X"07", X"8a", X"82", X"8e", X"83", X"8f", 
    X"f0", X"eb", X"12", X"66", X"a0", X"a3", X"ec", X"12", 
    X"66", X"a0", X"a3", X"ed", X"12", X"66", X"a0", X"d0", 
    X"07", X"d0", X"06", X"eb", X"4c", X"70", X"26", X"a8", 
    X"0c", X"08", X"86", X"03", X"08", X"86", X"04", X"08", 
    X"86", X"05", X"8b", X"82", X"8c", X"83", X"8d", X"f0", 
    X"c0", X"07", X"c0", X"06", X"12", X"62", X"2d", X"d0", 
    X"06", X"d0", X"07", X"a8", X"0c", X"08", X"e4", X"f6", 
    X"08", X"f6", X"08", X"76", X"00", X"a8", X"0c", X"08", 
    X"e6", X"08", X"46", X"70", X"03", X"02", X"03", X"b9", 
    X"e5", X"0c", X"24", X"f9", X"f8", X"86", X"02", X"08", 
    X"86", X"03", X"e4", X"fc", X"fd", X"c0", X"e0", X"c0", 
    X"e0", X"c0", X"e0", X"a8", X"0c", X"08", X"e6", X"c0", 
    X"e0", X"08", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"e5", X"0c", X"24", X"f2", X"f8", X"e6", X"c0", 
    X"e0", X"08", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"e5", X"0c", X"24", X"f5", X"f8", X"e6", X"c0", 
    X"e0", X"e5", X"0c", X"24", X"f6", X"f8", X"e6", X"c0", 
    X"e0", X"08", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"c0", X"02", X"c0", X"03", X"c0", X"04", X"c0", 
    X"05", X"e5", X"0c", X"24", X"fb", X"f8", X"e6", X"c0", 
    X"e0", X"08", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"8e", X"82", X"8f", X"83", X"12", X"03", X"c2", 
    X"e5", X"81", X"24", X"ec", X"f5", X"81", X"a8", X"0c", 
    X"08", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"06", X"bb", X"75", X"82", X"01", X"80", 
    X"03", X"75", X"82", X"ff", X"85", X"0c", X"81", X"d0", 
    X"0c", X"22", X"c0", X"0c", X"85", X"81", X"0c", X"c0", 
    X"82", X"c0", X"83", X"e5", X"81", X"24", X"0c", X"f5", 
    X"81", X"e5", X"0c", X"24", X"ed", X"f8", X"e5", X"0c", 
    X"24", X"09", X"f9", X"e6", X"f7", X"08", X"09", X"e6", 
    X"f7", X"08", X"09", X"e6", X"f7", X"e5", X"0c", X"24", 
    X"09", X"f8", X"74", X"20", X"26", X"fa", X"e4", X"08", 
    X"36", X"fe", X"08", X"86", X"07", X"8a", X"82", X"8e", 
    X"83", X"8f", X"f0", X"e5", X"0c", X"24", X"0c", X"f8", 
    X"12", X"70", X"5a", X"f6", X"a3", X"12", X"70", X"5a", 
    X"08", X"f6", X"a3", X"12", X"70", X"5a", X"08", X"f6", 
    X"e5", X"0c", X"24", X"0c", X"f8", X"e5", X"0c", X"24", 
    X"03", X"f9", X"e6", X"f7", X"08", X"09", X"e6", X"f7", 
    X"08", X"09", X"e6", X"f7", X"e5", X"0c", X"24", X"09", 
    X"f8", X"e5", X"0c", X"24", X"06", X"f9", X"74", X"2b", 
    X"26", X"f7", X"e4", X"08", X"36", X"09", X"f7", X"08", 
    X"09", X"e6", X"f7", X"e5", X"0c", X"24", X"f7", X"f8", 
    X"e6", X"24", X"ff", X"fa", X"08", X"e6", X"34", X"ff", 
    X"fe", X"08", X"e6", X"34", X"ff", X"08", X"e6", X"34", 
    X"ff", X"e5", X"0c", X"24", X"0c", X"f8", X"ea", X"26", 
    X"fa", X"ee", X"08", X"36", X"fe", X"08", X"86", X"05", 
    X"e5", X"0c", X"24", X"06", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"ea", X"12", X"66", 
    X"a0", X"a3", X"ee", X"12", X"66", X"a0", X"a3", X"ed", 
    X"12", X"66", X"a0", X"e5", X"0c", X"24", X"09", X"f8", 
    X"74", X"23", X"26", X"fd", X"e4", X"08", X"36", X"fe", 
    X"08", X"86", X"07", X"7b", X"00", X"e5", X"0c", X"24", 
    X"06", X"f8", X"eb", X"2d", X"f6", X"e4", X"3e", X"08", 
    X"f6", X"08", X"a6", X"07", X"c0", X"05", X"c0", X"06", 
    X"c0", X"07", X"e5", X"0c", X"24", X"fb", X"f8", X"eb", 
    X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", X"86", 
    X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"70", X"5a", X"fc", X"e5", X"0c", X"24", X"06", X"f8", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"ec", X"12", X"66", X"a0", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"70", X"5a", X"d0", X"07", X"d0", 
    X"06", X"d0", X"05", X"60", X"06", X"0b", X"bb", X"08", 
    X"00", X"40", X"aa", X"e5", X"0c", X"24", X"09", X"f8", 
    X"74", X"2a", X"26", X"fd", X"e4", X"08", X"36", X"fe", 
    X"08", X"86", X"07", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"e4", X"12", X"66", X"a0", X"e5", X"0c", X"24", 
    X"f3", X"f8", X"b6", X"04", X"00", X"40", X"07", X"e5", 
    X"0c", X"24", X"f3", X"f8", X"76", X"03", X"e5", X"0c", 
    X"24", X"09", X"f8", X"74", X"1f", X"26", X"fd", X"e4", 
    X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"e5", X"0c", X"24", X"f3", 
    X"f8", X"e6", X"12", X"66", X"a0", X"e5", X"0c", X"24", 
    X"09", X"f8", X"74", X"03", X"26", X"fd", X"e4", X"08", 
    X"36", X"fe", X"08", X"86", X"07", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"2c", X"bf", X"e5", X"0c", 
    X"24", X"09", X"f8", X"74", X"11", X"26", X"fd", X"e4", 
    X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"2c", X"bf", X"e5", 
    X"0c", X"24", X"09", X"f8", X"74", X"0b", X"26", X"fd", 
    X"e4", X"08", X"36", X"fe", X"08", X"86", X"07", X"e5", 
    X"0c", X"24", X"ed", X"f8", X"86", X"02", X"08", X"86", 
    X"03", X"08", X"86", X"04", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"ea", X"12", X"66", X"a0", X"a3", X"eb", 
    X"12", X"66", X"a0", X"a3", X"ec", X"12", X"66", X"a0", 
    X"e5", X"0c", X"24", X"09", X"f8", X"e5", X"0c", X"24", 
    X"06", X"f9", X"74", X"11", X"26", X"f7", X"e4", X"08", 
    X"36", X"09", X"f7", X"08", X"09", X"e6", X"f7", X"e5", 
    X"0c", X"24", X"f3", X"f8", X"86", X"07", X"7e", X"00", 
    X"74", X"04", X"c3", X"9f", X"ff", X"e4", X"9e", X"fe", 
    X"e5", X"0c", X"24", X"06", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"ef", X"12", X"66", 
    X"a0", X"a3", X"ee", X"12", X"66", X"a0", X"e5", X"0c", 
    X"24", X"09", X"f8", X"74", X"19", X"26", X"fd", X"e4", 
    X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"ea", X"12", X"66", X"a0", 
    X"a3", X"eb", X"12", X"66", X"a0", X"a3", X"ec", X"12", 
    X"66", X"a0", X"e5", X"0c", X"24", X"09", X"f8", X"74", 
    X"2e", X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", 
    X"86", X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"e4", X"12", X"66", X"a0", X"a3", X"12", X"66", X"a0", 
    X"a3", X"12", X"66", X"a0", X"a3", X"12", X"66", X"a0", 
    X"e5", X"0c", X"24", X"09", X"f8", X"74", X"32", X"26", 
    X"fd", X"e4", X"08", X"36", X"fe", X"08", X"86", X"07", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"e4", X"12", 
    X"66", X"a0", X"e5", X"0c", X"24", X"f4", X"f8", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"08", X"e6", 
    X"c0", X"e0", X"a8", X"0c", X"08", X"e6", X"c0", X"e0", 
    X"08", X"e6", X"c0", X"e0", X"e5", X"0c", X"24", X"03", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"62", X"4b", X"af", X"82", X"ae", X"83", 
    X"ad", X"f0", X"e5", X"81", X"24", X"fb", X"f5", X"81", 
    X"e5", X"0c", X"24", X"09", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"ef", X"12", X"66", 
    X"a0", X"a3", X"ee", X"12", X"66", X"a0", X"a3", X"ed", 
    X"12", X"66", X"a0", X"e5", X"0c", X"24", X"f0", X"f8", 
    X"e6", X"08", X"46", X"60", X"28", X"e5", X"0c", X"24", 
    X"f0", X"f8", X"86", X"05", X"08", X"86", X"06", X"08", 
    X"86", X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"e5", X"0c", X"24", X"09", X"f8", X"e6", X"12", X"66", 
    X"a0", X"a3", X"08", X"e6", X"12", X"66", X"a0", X"a3", 
    X"08", X"e6", X"12", X"66", X"a0", X"85", X"0c", X"81", 
    X"d0", X"0c", X"22", X"ad", X"82", X"ae", X"83", X"af", 
    X"f0", X"c0", X"e0", X"c0", X"a8", X"c2", X"af", X"90", 
    X"00", X"66", X"e0", X"24", X"01", X"f0", X"90", X"00", 
    X"09", X"e0", X"fa", X"a3", X"e0", X"fb", X"a3", X"e0", 
    X"fc", X"ea", X"4b", X"70", X"24", X"90", X"00", X"09", 
    X"ed", X"f0", X"ee", X"a3", X"f0", X"ef", X"a3", X"f0", 
    X"90", X"00", X"66", X"e0", X"fc", X"bc", X"01", X"55", 
    X"c0", X"07", X"c0", X"06", X"c0", X"05", X"12", X"14", 
    X"65", X"d0", X"05", X"d0", X"06", X"d0", X"07", X"80", 
    X"44", X"90", X"00", X"6a", X"e0", X"70", X"3e", X"90", 
    X"00", X"09", X"e0", X"fa", X"a3", X"e0", X"fb", X"a3", 
    X"e0", X"fc", X"74", X"1f", X"2a", X"fa", X"e4", X"3b", 
    X"fb", X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"12", 
    X"70", X"5a", X"fa", X"74", X"1f", X"2d", X"f9", X"e4", 
    X"3e", X"fb", X"8f", X"04", X"89", X"82", X"8b", X"83", 
    X"8c", X"f0", X"12", X"70", X"5a", X"f9", X"c3", X"9a", 
    X"40", X"0b", X"90", X"00", X"09", X"ed", X"f0", X"ee", 
    X"a3", X"f0", X"ef", X"a3", X"f0", X"90", X"00", X"6e", 
    X"e0", X"24", X"01", X"f0", X"74", X"1f", X"2d", X"fa", 
    X"e4", X"3e", X"fb", X"8f", X"04", X"8a", X"82", X"8b", 
    X"83", X"8c", X"f0", X"12", X"70", X"5a", X"f9", X"90", 
    X"00", X"69", X"e0", X"c3", X"99", X"50", X"05", X"90", 
    X"00", X"69", X"e9", X"f0", X"74", X"03", X"2d", X"fd", 
    X"e4", X"3e", X"fe", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"12", X"70", X"5a", X"75", X"f0", X"0c", X"a4", 
    X"24", X"0c", X"f8", X"74", X"00", X"35", X"f0", X"f9", 
    X"c0", X"02", X"c0", X"03", X"c0", X"04", X"7c", X"00", 
    X"c0", X"04", X"c0", X"03", X"c0", X"02", X"c0", X"05", 
    X"c0", X"06", X"c0", X"07", X"88", X"82", X"89", X"83", 
    X"8c", X"f0", X"12", X"2c", X"df", X"15", X"81", X"15", 
    X"81", X"15", X"81", X"d0", X"02", X"d0", X"03", X"d0", 
    X"04", X"d0", X"e0", X"53", X"e0", X"80", X"e5", X"e0", 
    X"42", X"a8", X"d0", X"e0", X"90", X"00", X"6a", X"e0", 
    X"d0", X"04", X"d0", X"03", X"d0", X"02", X"60", X"2e", 
    X"90", X"00", X"09", X"e0", X"fd", X"a3", X"e0", X"fe", 
    X"a3", X"e0", X"ff", X"74", X"1f", X"2d", X"fd", X"e4", 
    X"3e", X"fe", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"70", X"5a", X"fd", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"12", X"70", X"5a", X"fa", X"c3", X"ed", 
    X"9a", X"50", X"03", X"12", X"64", X"b5", X"22", X"c0", 
    X"0c", X"85", X"81", X"0c", X"c0", X"82", X"c0", X"83", 
    X"c0", X"f0", X"05", X"81", X"05", X"81", X"7e", X"00", 
    X"c0", X"06", X"12", X"09", X"4a", X"d0", X"06", X"90", 
    X"00", X"67", X"e0", X"fa", X"a3", X"e0", X"fb", X"e5", 
    X"0c", X"24", X"04", X"f8", X"a6", X"02", X"08", X"a6", 
    X"03", X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", X"fb", 
    X"a3", X"12", X"70", X"5a", X"fc", X"e5", X"0c", X"24", 
    X"fc", X"f8", X"e6", X"2b", X"fd", X"08", X"e6", X"3c", 
    X"ff", X"8d", X"02", X"e5", X"0c", X"24", X"04", X"f8", 
    X"c3", X"e6", X"9b", X"08", X"e6", X"9c", X"50", X"18", 
    X"c3", X"ea", X"9b", X"ef", X"9c", X"50", X"27", X"e5", 
    X"0c", X"24", X"04", X"f8", X"c3", X"e6", X"9a", X"08", 
    X"e6", X"9f", X"50", X"1a", X"7e", X"01", X"80", X"16", 
    X"c3", X"ea", X"9b", X"ef", X"9c", X"40", X"0d", X"e5", 
    X"0c", X"24", X"04", X"f8", X"c3", X"e6", X"9a", X"08", 
    X"e6", X"9f", X"50", X"02", X"7e", X"01", X"a8", X"0c", 
    X"08", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"ea", X"12", X"66", X"a0", X"a3", X"ef", X"12", 
    X"66", X"a0", X"ee", X"60", X"19", X"e5", X"0c", X"24", 
    X"04", X"f8", X"ea", X"c3", X"96", X"fa", X"ef", X"08", 
    X"96", X"ff", X"e4", X"c0", X"e0", X"8a", X"82", X"8f", 
    X"83", X"12", X"22", X"38", X"15", X"81", X"12", X"09", 
    X"52", X"e5", X"82", X"70", X"03", X"12", X"64", X"b5", 
    X"85", X"0c", X"81", X"d0", X"0c", X"22", X"ae", X"82", 
    X"af", X"83", X"7d", X"00", X"ee", X"4f", X"60", X"1e", 
    X"c0", X"07", X"c0", X"06", X"12", X"09", X"4a", X"d0", 
    X"06", X"d0", X"07", X"e4", X"c0", X"e0", X"8e", X"82", 
    X"8f", X"83", X"12", X"22", X"38", X"15", X"81", X"12", 
    X"09", X"52", X"af", X"82", X"8f", X"05", X"ed", X"70", 
    X"03", X"12", X"64", X"b5", X"22", X"74", X"71", X"c0", 
    X"e0", X"74", X"00", X"c0", X"e0", X"e4", X"c0", X"e0", 
    X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", 
    X"74", X"ba", X"c0", X"e0", X"e4", X"c0", X"e0", X"74", 
    X"eb", X"c0", X"e0", X"74", X"70", X"c0", X"e0", X"74", 
    X"80", X"c0", X"e0", X"90", X"14", X"54", X"12", X"02", 
    X"80", X"af", X"82", X"e5", X"81", X"24", X"f4", X"f5", 
    X"81", X"bf", X"01", X"1a", X"c2", X"af", X"90", X"00", 
    X"6f", X"74", X"ff", X"f0", X"a3", X"f0", X"90", X"00", 
    X"6a", X"74", X"01", X"f0", X"90", X"00", X"67", X"e4", 
    X"f0", X"a3", X"f0", X"12", X"64", X"41", X"22", X"c2", 
    X"af", X"90", X"00", X"6a", X"e4", X"f0", X"12", X"64", 
    X"b4", X"22", X"90", X"00", X"74", X"e0", X"24", X"01", 
    X"f0", X"22", X"c0", X"0c", X"e5", X"81", X"f5", X"0c", 
    X"24", X"06", X"f5", X"81", X"e5", X"0c", X"24", X"04", 
    X"f8", X"e4", X"f6", X"08", X"f6", X"08", X"76", X"00", 
    X"7c", X"00", X"c0", X"e0", X"c0", X"a8", X"c2", X"af", 
    X"90", X"00", X"74", X"e0", X"14", X"f0", X"e0", X"60", 
    X"03", X"02", X"0a", X"f7", X"90", X"00", X"66", X"e0", 
    X"70", X"03", X"02", X"0a", X"f7", X"90", X"00", X"5a", 
    X"e0", X"70", X"03", X"02", X"0a", X"b5", X"c0", X"04", 
    X"90", X"00", X"60", X"e0", X"fa", X"a3", X"e0", X"fb", 
    X"a3", X"e0", X"fc", X"74", X"08", X"2a", X"fa", X"e4", 
    X"3b", X"fb", X"8a", X"82", X"8b", X"83", X"8c", X"f0", 
    X"12", X"70", X"5a", X"fa", X"a3", X"12", X"70", X"5a", 
    X"fb", X"a3", X"12", X"70", X"5a", X"fc", X"e5", X"0c", 
    X"24", X"04", X"f8", X"a6", X"02", X"08", X"a6", X"03", 
    X"08", X"a6", X"04", X"e5", X"0c", X"24", X"04", X"f8", 
    X"74", X"11", X"26", X"fa", X"e4", X"08", X"36", X"fb", 
    X"08", X"86", X"04", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"c0", X"04", X"12", X"30", X"3b", X"d0", X"04", 
    X"e5", X"0c", X"24", X"04", X"f8", X"74", X"03", X"26", 
    X"fa", X"e4", X"08", X"36", X"fb", X"08", X"86", X"04", 
    X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"c0", X"04", 
    X"12", X"30", X"3b", X"d0", X"04", X"e5", X"0c", X"24", 
    X"04", X"f8", X"a9", X"0c", X"09", X"74", X"1f", X"26", 
    X"f7", X"e4", X"08", X"36", X"09", X"f7", X"08", X"09", 
    X"e6", X"f7", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"ff", X"90", X"00", X"69", X"e0", X"c3", X"9f", X"d0", 
    X"04", X"50", X"05", X"90", X"00", X"69", X"ef", X"f0", 
    X"c0", X"04", X"e5", X"0c", X"24", X"04", X"f8", X"74", 
    X"03", X"26", X"fa", X"e4", X"08", X"36", X"fb", X"08", 
    X"86", X"04", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"75", X"f0", X"0c", X"a4", X"24", X"0c", X"fe", X"74", 
    X"00", X"35", X"f0", X"ff", X"7d", X"00", X"c0", X"04", 
    X"c0", X"02", X"c0", X"03", X"c0", X"04", X"8e", X"82", 
    X"8f", X"83", X"8d", X"f0", X"12", X"2c", X"df", X"15", 
    X"81", X"15", X"81", X"15", X"81", X"d0", X"04", X"a8", 
    X"0c", X"08", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"12", X"70", X"5a", X"ff", X"90", X"00", 
    X"09", X"e0", X"fc", X"a3", X"e0", X"fd", X"a3", X"e0", 
    X"fe", X"74", X"1f", X"2c", X"fc", X"e4", X"3d", X"fd", 
    X"8c", X"82", X"8d", X"83", X"8e", X"f0", X"12", X"70", 
    X"5a", X"fc", X"c3", X"ef", X"9c", X"d0", X"04", X"50", 
    X"03", X"02", X"09", X"85", X"90", X"00", X"6c", X"74", 
    X"01", X"f0", X"02", X"09", X"85", X"e5", X"0c", X"24", 
    X"04", X"f8", X"e6", X"08", X"46", X"60", X"07", X"c0", 
    X"04", X"12", X"14", X"c0", X"d0", X"04", X"90", X"00", 
    X"6b", X"e0", X"ff", X"fe", X"60", X"1e", X"8e", X"07", 
    X"c0", X"07", X"c0", X"04", X"12", X"0b", X"66", X"e5", 
    X"82", X"d0", X"04", X"d0", X"07", X"60", X"06", X"90", 
    X"00", X"6c", X"74", X"01", X"f0", X"df", X"e9", X"90", 
    X"00", X"6b", X"e4", X"f0", X"90", X"00", X"6c", X"e0", 
    X"60", X"05", X"7c", X"01", X"12", X"64", X"b5", X"d0", 
    X"e0", X"53", X"e0", X"80", X"e5", X"e0", X"42", X"a8", 
    X"d0", X"e0", X"8c", X"82", X"85", X"0c", X"81", X"d0", 
    X"0c", X"22", X"c0", X"e0", X"c0", X"a8", X"c2", X"af", 
    X"90", X"00", X"67", X"e0", X"fe", X"a3", X"e0", X"ff", 
    X"d0", X"e0", X"53", X"e0", X"80", X"e5", X"e0", X"42", 
    X"a8", X"d0", X"e0", X"8e", X"82", X"8f", X"83", X"22", 
    X"90", X"00", X"67", X"e0", X"fe", X"a3", X"e0", X"8e", 
    X"82", X"f5", X"83", X"22", X"90", X"00", X"66", X"e0", 
    X"f5", X"82", X"22", X"ad", X"82", X"ae", X"83", X"af", 
    X"f0", X"ed", X"4e", X"70", X"0d", X"90", X"00", X"09", 
    X"e0", X"fa", X"a3", X"e0", X"fb", X"a3", X"e0", X"fc", 
    X"80", X"06", X"8d", X"02", X"8e", X"03", X"8f", X"04", 
    X"74", X"23", X"2a", X"fa", X"e4", X"3b", X"fb", X"8a", 
    X"82", X"8b", X"83", X"8c", X"f0", X"22", X"c0", X"0c", 
    X"e5", X"81", X"f5", X"0c", X"24", X"06", X"f5", X"81", 
    X"e5", X"0c", X"24", X"04", X"f8", X"76", X"00", X"90", 
    X"00", X"74", X"e0", X"60", X"03", X"02", X"0d", X"f2", 
    X"90", X"00", X"67", X"e0", X"fd", X"a3", X"e0", X"fe", 
    X"e5", X"0c", X"24", X"05", X"f8", X"74", X"01", X"2d", 
    X"f6", X"e4", X"3e", X"08", X"f6", X"e5", X"0c", X"24", 
    X"05", X"f8", X"90", X"00", X"67", X"e6", X"f0", X"08", 
    X"e6", X"a3", X"f0", X"e5", X"0c", X"24", X"05", X"f8", 
    X"e6", X"08", X"46", X"70", X"3a", X"90", X"00", X"54", 
    X"e0", X"fa", X"a3", X"e0", X"fb", X"a3", X"e0", X"fc", 
    X"8b", X"05", X"8c", X"06", X"90", X"00", X"57", X"e0", 
    X"fb", X"a3", X"e0", X"fc", X"a3", X"e0", X"ff", X"90", 
    X"00", X"54", X"eb", X"f0", X"ec", X"a3", X"f0", X"ef", 
    X"a3", X"f0", X"90", X"00", X"57", X"ea", X"f0", X"ed", 
    X"a3", X"f0", X"ee", X"a3", X"f0", X"90", X"00", X"6d", 
    X"e0", X"24", X"01", X"f0", X"12", X"14", X"c0", X"90", 
    X"00", X"6f", X"e0", X"fb", X"a3", X"e0", X"fc", X"e5", 
    X"0c", X"24", X"05", X"f8", X"c3", X"e6", X"9b", X"08", 
    X"e6", X"9c", X"50", X"03", X"02", X"0d", X"bb", X"90", 
    X"00", X"54", X"e0", X"fa", X"a3", X"e0", X"fb", X"a3", 
    X"e0", X"fc", X"8a", X"82", X"8b", X"83", X"8c", X"f0", 
    X"12", X"70", X"5a", X"70", X"0b", X"90", X"00", X"6f", 
    X"74", X"ff", X"f0", X"a3", X"f0", X"02", X"0d", X"bb", 
    X"90", X"00", X"54", X"e0", X"fa", X"a3", X"e0", X"fb", 
    X"a3", X"e0", X"fc", X"74", X"04", X"2a", X"fa", X"e4", 
    X"3b", X"fb", X"74", X"02", X"2a", X"fa", X"e4", X"3b", 
    X"fb", X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"12", 
    X"70", X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"fb", 
    X"a3", X"12", X"70", X"5a", X"fc", X"74", X"08", X"2a", 
    X"fa", X"e4", X"3b", X"fb", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"12", X"70", X"5a", X"fa", X"a3", X"12", 
    X"70", X"5a", X"fb", X"a3", X"12", X"70", X"5a", X"fc", 
    X"74", X"03", X"2a", X"fd", X"e4", X"3b", X"fe", X"8c", 
    X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"70", X"5a", X"ff", X"a3", X"12", X"70", X"5a", X"fe", 
    X"e5", X"0c", X"24", X"05", X"f8", X"c3", X"e6", X"9f", 
    X"08", X"e6", X"9e", X"50", X"0b", X"90", X"00", X"6f", 
    X"ef", X"f0", X"ee", X"a3", X"f0", X"02", X"0d", X"bb", 
    X"74", X"03", X"2a", X"fd", X"e4", X"3b", X"fe", X"8c", 
    X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"c0", 
    X"04", X"c0", X"03", X"c0", X"02", X"12", X"30", X"3b", 
    X"d0", X"02", X"d0", X"03", X"d0", X"04", X"a8", X"0c", 
    X"08", X"74", X"11", X"2a", X"f6", X"e4", X"3b", X"08", 
    X"f6", X"08", X"a6", X"04", X"74", X"1c", X"2a", X"fd", 
    X"e4", X"3b", X"fe", X"8c", X"07", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fd", X"a3", 
    X"12", X"70", X"5a", X"fe", X"a3", X"12", X"70", X"5a", 
    X"ed", X"4e", X"60", X"1a", X"a8", X"0c", X"08", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"c0", 
    X"04", X"c0", X"03", X"c0", X"02", X"12", X"30", X"3b", 
    X"d0", X"02", X"d0", X"03", X"d0", X"04", X"74", X"1f", 
    X"2a", X"fd", X"e4", X"3b", X"fe", X"8c", X"07", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"a8", X"0c", X"08", 
    X"12", X"70", X"5a", X"f6", X"c0", X"02", X"c0", X"03", 
    X"c0", X"04", X"90", X"00", X"69", X"e0", X"fc", X"a8", 
    X"0c", X"08", X"c3", X"ec", X"96", X"d0", X"04", X"d0", 
    X"03", X"d0", X"02", X"50", X"08", X"a8", X"0c", X"08", 
    X"90", X"00", X"69", X"e6", X"f0", X"a8", X"0c", X"08", 
    X"74", X"03", X"2a", X"f6", X"e4", X"3b", X"08", X"f6", 
    X"08", X"a6", X"04", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"12", X"70", X"5a", X"75", X"f0", X"0c", X"a4", 
    X"24", X"0c", X"fb", X"74", X"00", X"35", X"f0", X"fc", 
    X"7a", X"00", X"c0", X"07", X"c0", X"06", X"c0", X"05", 
    X"a8", X"0c", X"08", X"e6", X"c0", X"e0", X"08", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"8b", X"82", 
    X"8c", X"83", X"8a", X"f0", X"12", X"2c", X"df", X"15", 
    X"81", X"15", X"81", X"15", X"81", X"d0", X"05", X"d0", 
    X"06", X"d0", X"07", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"12", X"70", X"5a", X"fd", X"90", X"00", X"09", 
    X"e0", X"fc", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", 
    X"74", X"1f", X"2c", X"fc", X"e4", X"3e", X"fe", X"8c", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"fc", X"c3", X"ed", X"9c", X"50", X"03", X"02", X"0b", 
    X"ff", X"e5", X"0c", X"24", X"04", X"f8", X"76", X"01", 
    X"02", X"0b", X"ff", X"90", X"00", X"09", X"e0", X"fd", 
    X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"74", X"1f", 
    X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"70", X"5a", X"75", X"f0", 
    X"0c", X"a4", X"24", X"0c", X"f5", X"82", X"74", X"00", 
    X"35", X"f0", X"f5", X"83", X"e0", X"24", X"fe", X"50", 
    X"10", X"e5", X"0c", X"24", X"04", X"f8", X"76", X"01", 
    X"80", X"07", X"90", X"00", X"6b", X"e0", X"24", X"01", 
    X"f0", X"90", X"00", X"6c", X"e0", X"60", X"07", X"e5", 
    X"0c", X"24", X"04", X"f8", X"76", X"01", X"e5", X"0c", 
    X"24", X"04", X"f8", X"86", X"82", X"85", X"0c", X"81", 
    X"d0", X"0c", X"22", X"c0", X"0c", X"e5", X"81", X"f5", 
    X"0c", X"24", X"0a", X"f5", X"81", X"90", X"00", X"74", 
    X"e0", X"60", X"09", X"90", X"00", X"6c", X"74", X"01", 
    X"f0", X"02", X"0f", X"8c", X"90", X"00", X"6c", X"e4", 
    X"f0", X"90", X"00", X"69", X"e0", X"ff", X"ef", X"75", 
    X"f0", X"0c", X"a4", X"fd", X"ae", X"f0", X"24", X"0c", 
    X"fb", X"ee", X"34", X"00", X"fc", X"8b", X"82", X"8c", 
    X"83", X"e0", X"70", X"03", X"1f", X"80", X"e7", X"e5", 
    X"0c", X"24", X"07", X"f8", X"a6", X"07", X"ed", X"24", 
    X"0c", X"fd", X"ee", X"34", X"00", X"fe", X"e5", X"0c", 
    X"24", X"08", X"f8", X"a6", X"05", X"08", X"a6", X"06", 
    X"08", X"76", X"00", X"e5", X"0c", X"24", X"08", X"f8", 
    X"74", X"01", X"26", X"fa", X"e4", X"08", X"36", X"fb", 
    X"08", X"86", X"07", X"8a", X"82", X"8b", X"83", X"8f", 
    X"f0", X"12", X"70", X"5a", X"fc", X"a3", X"12", X"70", 
    X"5a", X"fd", X"a3", X"12", X"70", X"5a", X"fe", X"74", 
    X"02", X"2c", X"fc", X"e4", X"3d", X"fd", X"8c", X"82", 
    X"8d", X"83", X"8e", X"f0", X"12", X"70", X"5a", X"fc", 
    X"a3", X"12", X"70", X"5a", X"fd", X"a3", X"12", X"70", 
    X"5a", X"fe", X"8a", X"82", X"8b", X"83", X"8f", X"f0", 
    X"ec", X"12", X"66", X"a0", X"a3", X"ed", X"12", X"66", 
    X"a0", X"a3", X"ee", X"12", X"66", X"a0", X"8a", X"82", 
    X"8b", X"83", X"8f", X"f0", X"a8", X"0c", X"08", X"12", 
    X"70", X"5a", X"f6", X"a3", X"12", X"70", X"5a", X"08", 
    X"f6", X"a3", X"12", X"70", X"5a", X"08", X"f6", X"e5", 
    X"0c", X"24", X"04", X"f8", X"a6", X"04", X"08", X"a6", 
    X"05", X"08", X"a6", X"06", X"e5", X"0c", X"24", X"08", 
    X"f8", X"74", X"04", X"26", X"fc", X"e4", X"08", X"36", 
    X"fd", X"08", X"86", X"06", X"e5", X"0c", X"24", X"04", 
    X"f8", X"c0", X"04", X"c0", X"05", X"c0", X"06", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"12", 
    X"00", X"11", X"15", X"81", X"15", X"81", X"15", X"81", 
    X"70", X"36", X"a8", X"0c", X"08", X"74", X"02", X"26", 
    X"fc", X"e4", X"08", X"36", X"fd", X"08", X"86", X"06", 
    X"8c", X"82", X"8d", X"83", X"8e", X"f0", X"12", X"70", 
    X"5a", X"fc", X"a3", X"12", X"70", X"5a", X"fd", X"a3", 
    X"12", X"70", X"5a", X"fe", X"8a", X"82", X"8b", X"83", 
    X"8f", X"f0", X"ec", X"12", X"66", X"a0", X"a3", X"ed", 
    X"12", X"66", X"a0", X"a3", X"ee", X"12", X"66", X"a0", 
    X"8a", X"82", X"8b", X"83", X"8f", X"f0", X"12", X"70", 
    X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"fb", X"a3", 
    X"12", X"70", X"5a", X"ff", X"74", X"08", X"2a", X"fa", 
    X"e4", X"3b", X"fb", X"8a", X"82", X"8b", X"83", X"8f", 
    X"f0", X"12", X"70", X"5a", X"fa", X"a3", X"12", X"70", 
    X"5a", X"fb", X"a3", X"12", X"70", X"5a", X"ff", X"90", 
    X"00", X"09", X"ea", X"f0", X"eb", X"a3", X"f0", X"ef", 
    X"a3", X"f0", X"e5", X"0c", X"24", X"07", X"f8", X"90", 
    X"00", X"69", X"e6", X"f0", X"85", X"0c", X"81", X"d0", 
    X"0c", X"22", X"c0", X"0c", X"85", X"81", X"0c", X"ad", 
    X"82", X"ae", X"83", X"af", X"f0", X"90", X"00", X"09", 
    X"e0", X"fa", X"a3", X"e0", X"fb", X"a3", X"e0", X"fc", 
    X"74", X"11", X"2a", X"fa", X"e4", X"3b", X"fb", X"c0", 
    X"02", X"c0", X"03", X"c0", X"04", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"2e", X"3d", X"15", X"81", 
    X"15", X"81", X"15", X"81", X"74", X"01", X"c0", X"e0", 
    X"e5", X"0c", X"24", X"fc", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"12", X"22", X"38", X"15", X"81", X"d0", 
    X"0c", X"22", X"c0", X"0c", X"85", X"81", X"0c", X"c0", 
    X"82", X"c0", X"83", X"c0", X"f0", X"90", X"00", X"09", 
    X"e0", X"fa", X"a3", X"e0", X"fb", X"a3", X"e0", X"fc", 
    X"74", X"11", X"2a", X"fa", X"e4", X"3b", X"fb", X"e5", 
    X"0c", X"24", X"fc", X"f8", X"86", X"06", X"74", X"80", 
    X"08", X"46", X"ff", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"ee", X"12", X"66", X"a0", X"a3", X"ef", X"12", 
    X"66", X"a0", X"90", X"00", X"09", X"e0", X"fd", X"a3", 
    X"e0", X"fe", X"a3", X"e0", X"ff", X"74", X"11", X"2d", 
    X"fd", X"e4", X"3e", X"fe", X"c0", X"05", X"c0", X"06", 
    X"c0", X"07", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"2c", X"df", 
    X"15", X"81", X"15", X"81", X"15", X"81", X"74", X"01", 
    X"c0", X"e0", X"e5", X"0c", X"24", X"fa", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"12", X"22", X"38", X"15", 
    X"81", X"85", X"0c", X"81", X"d0", X"0c", X"22", X"c0", 
    X"0c", X"85", X"81", X"0c", X"05", X"81", X"05", X"81", 
    X"05", X"81", X"ad", X"82", X"ae", X"83", X"af", X"f0", 
    X"74", X"04", X"2d", X"fd", X"e4", X"3e", X"fe", X"74", 
    X"02", X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fd", 
    X"a3", X"12", X"70", X"5a", X"fe", X"a3", X"12", X"70", 
    X"5a", X"ff", X"74", X"08", X"2d", X"fd", X"e4", X"3e", 
    X"fe", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"70", X"5a", X"fd", X"a3", X"12", X"70", X"5a", X"fe", 
    X"a3", X"12", X"70", X"5a", X"ff", X"a8", X"0c", X"08", 
    X"a6", X"05", X"08", X"a6", X"06", X"08", X"a6", X"07", 
    X"a8", X"0c", X"08", X"74", X"11", X"26", X"fa", X"e4", 
    X"08", X"36", X"fb", X"08", X"86", X"04", X"8a", X"82", 
    X"8b", X"83", X"8c", X"f0", X"12", X"30", X"3b", X"90", 
    X"00", X"74", X"e0", X"60", X"03", X"02", X"11", X"48", 
    X"a8", X"0c", X"08", X"74", X"03", X"26", X"fa", X"e4", 
    X"08", X"36", X"fb", X"08", X"86", X"04", X"8a", X"82", 
    X"8b", X"83", X"8c", X"f0", X"12", X"30", X"3b", X"a8", 
    X"0c", X"08", X"74", X"1f", X"26", X"fa", X"e4", X"08", 
    X"36", X"fb", X"08", X"86", X"04", X"8a", X"82", X"8b", 
    X"83", X"8c", X"f0", X"12", X"70", X"5a", X"fe", X"90", 
    X"00", X"69", X"e0", X"c3", X"9e", X"50", X"05", X"90", 
    X"00", X"69", X"ee", X"f0", X"a8", X"0c", X"08", X"74", 
    X"03", X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", 
    X"86", X"07", X"8a", X"82", X"8b", X"83", X"8c", X"f0", 
    X"12", X"70", X"5a", X"75", X"f0", X"0c", X"a4", X"24", 
    X"0c", X"fb", X"74", X"00", X"35", X"f0", X"fc", X"7a", 
    X"00", X"c0", X"05", X"c0", X"06", X"c0", X"07", X"8b", 
    X"82", X"8c", X"83", X"8a", X"f0", X"12", X"2c", X"df", 
    X"15", X"81", X"15", X"81", X"15", X"81", X"80", X"23", 
    X"a8", X"0c", X"08", X"74", X"11", X"26", X"fd", X"e4", 
    X"08", X"36", X"fe", X"08", X"86", X"07", X"c0", X"05", 
    X"c0", X"06", X"c0", X"07", X"90", X"00", X"5a", X"75", 
    X"f0", X"00", X"12", X"2c", X"df", X"15", X"81", X"15", 
    X"81", X"15", X"81", X"a8", X"0c", X"08", X"74", X"1f", 
    X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", X"86", 
    X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"70", X"5a", X"fd", X"90", X"00", X"09", X"e0", X"fc", 
    X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"74", X"1f", 
    X"2c", X"fc", X"e4", X"3e", X"fe", X"8c", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"70", X"5a", X"c3", X"9d", 
    X"50", X"09", X"7f", X"01", X"90", X"00", X"6c", X"ef", 
    X"f0", X"80", X"02", X"7f", X"00", X"8f", X"82", X"85", 
    X"0c", X"81", X"d0", X"0c", X"22", X"c0", X"0c", X"e5", 
    X"81", X"f5", X"0c", X"24", X"06", X"f5", X"81", X"ad", 
    X"82", X"ae", X"83", X"af", X"f0", X"e5", X"0c", X"24", 
    X"fc", X"f8", X"86", X"03", X"74", X"80", X"08", X"46", 
    X"fc", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"eb", 
    X"12", X"66", X"a0", X"a3", X"ec", X"12", X"66", X"a0", 
    X"74", X"08", X"2d", X"fa", X"e4", X"3e", X"fb", X"8f", 
    X"04", X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"12", 
    X"70", X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"fb", 
    X"a3", X"12", X"70", X"5a", X"fc", X"e5", X"0c", X"24", 
    X"04", X"f8", X"a6", X"02", X"08", X"a6", X"03", X"08", 
    X"a6", X"04", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"30", X"3b", X"e5", X"0c", X"24", X"04", X"f8", 
    X"74", X"03", X"26", X"fd", X"e4", X"08", X"36", X"fe", 
    X"08", X"86", X"07", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"12", X"30", X"3b", X"e5", X"0c", X"24", X"04", 
    X"f8", X"74", X"1f", X"26", X"fd", X"e4", X"08", X"36", 
    X"fe", X"08", X"86", X"07", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"70", X"5a", X"fb", X"90", X"00", 
    X"69", X"e0", X"c3", X"9b", X"50", X"05", X"90", X"00", 
    X"69", X"eb", X"f0", X"e5", X"0c", X"24", X"04", X"f8", 
    X"a9", X"0c", X"09", X"74", X"03", X"26", X"f7", X"e4", 
    X"08", X"36", X"09", X"f7", X"08", X"09", X"e6", X"f7", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", 
    X"5a", X"75", X"f0", X"0c", X"a4", X"24", X"0c", X"fb", 
    X"74", X"00", X"35", X"f0", X"fc", X"7a", X"00", X"c0", 
    X"07", X"c0", X"06", X"c0", X"05", X"a8", X"0c", X"08", 
    X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"8b", X"82", X"8c", X"83", X"8a", 
    X"f0", X"12", X"2c", X"df", X"15", X"81", X"15", X"81", 
    X"15", X"81", X"d0", X"05", X"d0", X"06", X"d0", X"07", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", 
    X"5a", X"fd", X"90", X"00", X"09", X"e0", X"fc", X"a3", 
    X"e0", X"fe", X"a3", X"e0", X"ff", X"74", X"1f", X"2c", 
    X"fc", X"e4", X"3e", X"fe", X"8c", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"70", X"5a", X"c3", X"9d", X"50", 
    X"06", X"90", X"00", X"6c", X"74", X"01", X"f0", X"85", 
    X"0c", X"81", X"d0", X"0c", X"22", X"ad", X"82", X"ae", 
    X"83", X"af", X"f0", X"c0", X"e0", X"c0", X"a8", X"c2", 
    X"af", X"90", X"00", X"6d", X"e0", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"66", X"a0", X"0d", X"bd", 
    X"00", X"01", X"0e", X"90", X"00", X"67", X"e0", X"fb", 
    X"a3", X"e0", X"fc", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"eb", X"12", X"66", X"a0", X"a3", X"ec", X"12", 
    X"66", X"a0", X"d0", X"e0", X"53", X"e0", X"80", X"e5", 
    X"e0", X"42", X"a8", X"d0", X"e0", X"22", X"ad", X"82", 
    X"ae", X"83", X"af", X"f0", X"90", X"00", X"6d", X"e0", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"66", 
    X"a0", X"0d", X"bd", X"00", X"01", X"0e", X"90", X"00", 
    X"67", X"e0", X"fb", X"a3", X"e0", X"fc", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"eb", X"12", X"66", X"a0", 
    X"a3", X"ec", X"12", X"66", X"a0", X"22", X"c0", X"0c", 
    X"85", X"81", X"0c", X"c0", X"82", X"c0", X"83", X"c0", 
    X"f0", X"e5", X"81", X"24", X"04", X"f5", X"81", X"c0", 
    X"e0", X"c0", X"a8", X"c2", X"af", X"90", X"00", X"67", 
    X"e0", X"fb", X"a3", X"e0", X"fc", X"e5", X"0c", X"24", 
    X"06", X"f8", X"a6", X"03", X"08", X"a6", X"04", X"a8", 
    X"0c", X"08", X"74", X"01", X"26", X"fb", X"e4", X"08", 
    X"36", X"fa", X"08", X"86", X"04", X"8b", X"82", X"8a", 
    X"83", X"8c", X"f0", X"12", X"70", X"5a", X"fb", X"a3", 
    X"12", X"70", X"5a", X"fc", X"e5", X"0c", X"24", X"06", 
    X"f8", X"e6", X"c3", X"9b", X"fe", X"08", X"e6", X"9c", 
    X"ff", X"8e", X"02", X"a8", X"0c", X"08", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"70", 
    X"5a", X"fe", X"90", X"00", X"6d", X"e0", X"fd", X"b5", 
    X"06", X"02", X"80", X"11", X"e5", X"0c", X"24", X"06", 
    X"f8", X"c3", X"e6", X"9b", X"08", X"e6", X"9c", X"40", 
    X"04", X"7e", X"01", X"80", X"6d", X"e5", X"0c", X"24", 
    X"fb", X"f8", X"86", X"03", X"08", X"86", X"04", X"08", 
    X"86", X"05", X"8b", X"82", X"8c", X"83", X"8d", X"f0", 
    X"e5", X"0c", X"24", X"04", X"f8", X"12", X"70", X"5a", 
    X"f6", X"a3", X"12", X"70", X"5a", X"08", X"f6", X"e5", 
    X"0c", X"24", X"04", X"f8", X"c3", X"ea", X"96", X"ef", 
    X"08", X"96", X"50", X"2e", X"e5", X"0c", X"24", X"04", 
    X"f8", X"e6", X"c3", X"9a", X"fa", X"08", X"e6", X"9f", 
    X"ff", X"8b", X"82", X"8c", X"83", X"8d", X"f0", X"ea", 
    X"12", X"66", X"a0", X"a3", X"ef", X"12", X"66", X"a0", 
    X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"13", X"1e", X"7e", X"00", 
    X"80", X"10", X"8b", X"82", X"8c", X"83", X"8d", X"f0", 
    X"e4", X"12", X"66", X"a0", X"a3", X"12", X"66", X"a0", 
    X"7e", X"01", X"d0", X"e0", X"53", X"e0", X"80", X"e5", 
    X"e0", X"42", X"a8", X"d0", X"e0", X"8e", X"82", X"85", 
    X"0c", X"81", X"d0", X"0c", X"22", X"90", X"00", X"6c", 
    X"74", X"01", X"f0", X"22", X"12", X"14", X"bf", X"90", 
    X"00", X"0c", X"e0", X"24", X"fe", X"50", X"f5", X"12", 
    X"64", X"b5", X"80", X"f0", X"22", X"7f", X"00", X"ef", 
    X"75", X"f0", X"0c", X"a4", X"24", X"0c", X"fd", X"74", 
    X"00", X"35", X"f0", X"fe", X"7c", X"00", X"8d", X"82", 
    X"8e", X"83", X"8c", X"f0", X"c0", X"07", X"12", X"2b", 
    X"dd", X"d0", X"07", X"0f", X"bf", X"04", X"00", X"40", 
    X"de", X"90", X"00", X"3c", X"75", X"f0", X"00", X"12", 
    X"2b", X"dd", X"90", X"00", X"48", X"75", X"f0", X"00", 
    X"12", X"2b", X"dd", X"90", X"00", X"5a", X"75", X"f0", 
    X"00", X"12", X"2b", X"dd", X"90", X"00", X"54", X"74", 
    X"3c", X"f0", X"74", X"00", X"a3", X"f0", X"e4", X"a3", 
    X"f0", X"90", X"00", X"57", X"74", X"48", X"f0", X"74", 
    X"00", X"a3", X"f0", X"e4", X"a3", X"f0", X"22", X"22", 
    X"90", X"00", X"54", X"e0", X"fd", X"a3", X"e0", X"fe", 
    X"a3", X"e0", X"ff", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"12", X"70", X"5a", X"70", X"0a", X"90", X"00", 
    X"6f", X"74", X"ff", X"f0", X"a3", X"f0", X"80", X"66", 
    X"90", X"00", X"54", X"e0", X"fd", X"a3", X"e0", X"fe", 
    X"a3", X"e0", X"ff", X"74", X"04", X"2d", X"fd", X"e4", 
    X"3e", X"fe", X"74", X"02", X"2d", X"fd", X"e4", X"3e", 
    X"fe", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"70", X"5a", X"fd", X"a3", X"12", X"70", X"5a", X"fe", 
    X"a3", X"12", X"70", X"5a", X"ff", X"74", X"08", X"2d", 
    X"fd", X"e4", X"3e", X"fe", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"70", X"5a", X"fd", X"a3", X"12", 
    X"70", X"5a", X"fe", X"a3", X"12", X"70", X"5a", X"ff", 
    X"74", X"03", X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"fd", X"a3", X"12", X"70", X"5a", X"fe", X"90", X"00", 
    X"6f", X"ed", X"f0", X"ee", X"a3", X"f0", X"22", X"90", 
    X"00", X"09", X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", 
    X"e0", X"ff", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"22", X"c0", X"0c", X"85", X"81", X"0c", X"05", X"81", 
    X"05", X"81", X"90", X"00", X"09", X"e0", X"fd", X"a3", 
    X"e0", X"fe", X"a3", X"e0", X"ff", X"74", X"11", X"2d", 
    X"fd", X"e4", X"3e", X"fe", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"a8", X"0c", X"08", X"12", X"70", X"5a", 
    X"f6", X"a3", X"12", X"70", X"5a", X"08", X"f6", X"90", 
    X"00", X"09", X"e0", X"fb", X"a3", X"e0", X"fc", X"a3", 
    X"e0", X"ff", X"74", X"11", X"2b", X"fb", X"e4", X"3c", 
    X"fc", X"90", X"00", X"09", X"e0", X"fa", X"a3", X"e0", 
    X"fd", X"a3", X"e0", X"fe", X"74", X"1f", X"2a", X"fa", 
    X"e4", X"3d", X"fd", X"8a", X"82", X"8d", X"83", X"8e", 
    X"f0", X"12", X"70", X"5a", X"fa", X"7e", X"00", X"74", 
    X"04", X"c3", X"9a", X"fa", X"e4", X"9e", X"fe", X"8b", 
    X"82", X"8c", X"83", X"8f", X"f0", X"ea", X"12", X"66", 
    X"a0", X"a3", X"ee", X"12", X"66", X"a0", X"a8", X"0c", 
    X"08", X"86", X"82", X"08", X"86", X"83", X"85", X"0c", 
    X"81", X"d0", X"0c", X"22", X"c0", X"0c", X"e5", X"81", 
    X"f5", X"0c", X"24", X"07", X"f5", X"81", X"af", X"82", 
    X"c0", X"e0", X"c0", X"a8", X"c2", X"af", X"90", X"00", 
    X"09", X"e0", X"fc", X"a3", X"e0", X"fd", X"a3", X"e0", 
    X"fe", X"74", X"2e", X"2c", X"fc", X"e4", X"3d", X"fd", 
    X"8c", X"82", X"8d", X"83", X"8e", X"f0", X"12", X"70", 
    X"5a", X"fc", X"a3", X"12", X"70", X"5a", X"fd", X"a3", 
    X"12", X"70", X"5a", X"fe", X"a3", X"12", X"70", X"5a", 
    X"fb", X"ec", X"4d", X"4e", X"4b", X"70", X"41", X"90", 
    X"00", X"09", X"e0", X"fc", X"a3", X"e0", X"fd", X"a3", 
    X"e0", X"fe", X"74", X"32", X"2c", X"fc", X"e4", X"3d", 
    X"fd", X"8c", X"82", X"8d", X"83", X"8e", X"f0", X"74", 
    X"01", X"12", X"66", X"a0", X"e5", X"0c", X"24", X"fc", 
    X"f8", X"e6", X"08", X"46", X"60", X"1a", X"c0", X"07", 
    X"74", X"01", X"c0", X"e0", X"e5", X"0c", X"24", X"fc", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"12", X"22", 
    X"38", X"15", X"81", X"d0", X"07", X"12", X"64", X"b5", 
    X"d0", X"e0", X"53", X"e0", X"80", X"e5", X"e0", X"42", 
    X"a8", X"d0", X"e0", X"c0", X"e0", X"c0", X"a8", X"c2", 
    X"af", X"90", X"00", X"09", X"e0", X"fe", X"a3", X"e0", 
    X"fc", X"a3", X"e0", X"fd", X"74", X"2e", X"2e", X"fe", 
    X"e4", X"3c", X"fc", X"8e", X"82", X"8c", X"83", X"8d", 
    X"f0", X"e5", X"0c", X"24", X"04", X"f8", X"12", X"70", 
    X"5a", X"f6", X"a3", X"12", X"70", X"5a", X"08", X"f6", 
    X"a3", X"12", X"70", X"5a", X"08", X"f6", X"a3", X"12", 
    X"70", X"5a", X"08", X"f6", X"e5", X"0c", X"24", X"04", 
    X"f8", X"e6", X"08", X"46", X"08", X"46", X"08", X"46", 
    X"70", X"03", X"02", X"17", X"31", X"ef", X"60", X"2a", 
    X"90", X"00", X"09", X"e0", X"fa", X"a3", X"e0", X"fe", 
    X"a3", X"e0", X"ff", X"74", X"2e", X"2a", X"fa", X"e4", 
    X"3e", X"fe", X"8a", X"82", X"8e", X"83", X"8f", X"f0", 
    X"e4", X"12", X"66", X"a0", X"a3", X"12", X"66", X"a0", 
    X"a3", X"12", X"66", X"a0", X"a3", X"12", X"66", X"a0", 
    X"80", X"4f", X"90", X"00", X"09", X"e0", X"fa", X"a3", 
    X"e0", X"fe", X"a3", X"e0", X"ff", X"a8", X"0c", X"08", 
    X"74", X"2e", X"2a", X"f6", X"e4", X"3e", X"08", X"f6", 
    X"08", X"a6", X"07", X"e5", X"0c", X"24", X"04", X"f8", 
    X"e6", X"24", X"ff", X"fb", X"08", X"e6", X"34", X"ff", 
    X"fc", X"08", X"e6", X"34", X"ff", X"fd", X"08", X"e6", 
    X"34", X"ff", X"ff", X"a8", X"0c", X"08", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"eb", X"12", 
    X"66", X"a0", X"a3", X"ec", X"12", X"66", X"a0", X"a3", 
    X"ed", X"12", X"66", X"a0", X"a3", X"ef", X"12", X"66", 
    X"a0", X"90", X"00", X"09", X"e0", X"fd", X"a3", X"e0", 
    X"fe", X"a3", X"e0", X"ff", X"74", X"32", X"2d", X"fd", 
    X"e4", X"3e", X"fe", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"e4", X"12", X"66", X"a0", X"d0", X"e0", X"53", 
    X"e0", X"80", X"e5", X"e0", X"42", X"a8", X"d0", X"e0", 
    X"e5", X"0c", X"24", X"04", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"08", X"e6", X"85", 
    X"0c", X"81", X"d0", X"0c", X"22", X"c0", X"0c", X"85", 
    X"81", X"0c", X"c0", X"82", X"c0", X"83", X"c0", X"f0", 
    X"c0", X"e0", X"e5", X"81", X"24", X"0b", X"f5", X"81", 
    X"c0", X"e0", X"c0", X"a8", X"c2", X"af", X"90", X"00", 
    X"09", X"e0", X"fa", X"a3", X"e0", X"fb", X"a3", X"e0", 
    X"ff", X"74", X"32", X"2a", X"fa", X"e4", X"3b", X"fb", 
    X"8a", X"82", X"8b", X"83", X"8f", X"f0", X"12", X"70", 
    X"5a", X"fa", X"ba", X"02", X"03", X"02", X"18", X"79", 
    X"90", X"00", X"09", X"e0", X"fd", X"a3", X"e0", X"fe", 
    X"a3", X"e0", X"ff", X"e5", X"0c", X"24", X"05", X"f8", 
    X"74", X"2e", X"2d", X"f6", X"e4", X"3e", X"08", X"f6", 
    X"08", X"a6", X"07", X"90", X"00", X"09", X"e0", X"fa", 
    X"a3", X"e0", X"fb", X"a3", X"e0", X"fc", X"74", X"2e", 
    X"2a", X"fa", X"e4", X"3b", X"fb", X"8a", X"82", X"8b", 
    X"83", X"8c", X"f0", X"e5", X"0c", X"24", X"08", X"f8", 
    X"12", X"70", X"5a", X"f6", X"a3", X"12", X"70", X"5a", 
    X"08", X"f6", X"a3", X"12", X"70", X"5a", X"08", X"f6", 
    X"a3", X"12", X"70", X"5a", X"08", X"f6", X"a8", X"0c", 
    X"08", X"e6", X"f4", X"fd", X"08", X"e6", X"f4", X"fe", 
    X"08", X"e6", X"f4", X"fc", X"08", X"e6", X"f4", X"ff", 
    X"e5", X"0c", X"24", X"08", X"f8", X"e6", X"52", X"05", 
    X"08", X"e6", X"52", X"06", X"08", X"e6", X"52", X"04", 
    X"08", X"e6", X"52", X"07", X"e5", X"0c", X"24", X"05", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"ed", X"12", X"66", X"a0", X"a3", X"ee", X"12", 
    X"66", X"a0", X"a3", X"ec", X"12", X"66", X"a0", X"a3", 
    X"ef", X"12", X"66", X"a0", X"90", X"00", X"09", X"e0", 
    X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"74", 
    X"32", X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"74", X"01", X"12", X"66", 
    X"a0", X"e5", X"0c", X"24", X"f5", X"f8", X"e6", X"08", 
    X"46", X"60", X"16", X"74", X"01", X"c0", X"e0", X"e5", 
    X"0c", X"24", X"f5", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"12", X"22", X"38", X"15", X"81", X"12", X"64", 
    X"b5", X"d0", X"e0", X"53", X"e0", X"80", X"e5", X"e0", 
    X"42", X"a8", X"d0", X"e0", X"c0", X"e0", X"c0", X"a8", 
    X"c2", X"af", X"e5", X"0c", X"24", X"f7", X"f8", X"e6", 
    X"08", X"46", X"60", X"5f", X"e5", X"0c", X"24", X"f7", 
    X"f8", X"e5", X"0c", X"24", X"08", X"f9", X"e6", X"f7", 
    X"08", X"09", X"e6", X"f7", X"08", X"09", X"e6", X"f7", 
    X"90", X"00", X"09", X"e0", X"fa", X"a3", X"e0", X"fb", 
    X"a3", X"e0", X"fc", X"74", X"2e", X"2a", X"fa", X"e4", 
    X"3b", X"fb", X"8a", X"82", X"8b", X"83", X"8c", X"f0", 
    X"12", X"70", X"5a", X"fa", X"a3", X"12", X"70", X"5a", 
    X"fb", X"a3", X"12", X"70", X"5a", X"fc", X"a3", X"12", 
    X"70", X"5a", X"ff", X"e5", X"0c", X"24", X"08", X"f8", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"ea", X"12", X"66", X"a0", X"a3", X"eb", X"12", X"66", 
    X"a0", X"a3", X"ec", X"12", X"66", X"a0", X"a3", X"ef", 
    X"12", X"66", X"a0", X"90", X"00", X"09", X"e0", X"fd", 
    X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"74", X"32", 
    X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fd", X"bd", 
    X"02", X"02", X"80", X"05", X"7f", X"00", X"02", X"19", 
    X"b1", X"90", X"00", X"09", X"e0", X"fc", X"a3", X"e0", 
    X"fd", X"a3", X"e0", X"fe", X"e5", X"0c", X"24", X"08", 
    X"f8", X"74", X"2e", X"2c", X"f6", X"e4", X"3d", X"08", 
    X"f6", X"08", X"a6", X"06", X"90", X"00", X"09", X"e0", 
    X"fa", X"a3", X"e0", X"fb", X"a3", X"e0", X"fe", X"74", 
    X"2e", X"2a", X"fa", X"e4", X"3b", X"fb", X"8a", X"82", 
    X"8b", X"83", X"8e", X"f0", X"e5", X"0c", X"24", X"0c", 
    X"f8", X"12", X"70", X"5a", X"f6", X"a3", X"12", X"70", 
    X"5a", X"08", X"f6", X"a3", X"12", X"70", X"5a", X"08", 
    X"f6", X"a3", X"12", X"70", X"5a", X"08", X"f6", X"e5", 
    X"0c", X"24", X"fa", X"f8", X"e6", X"f4", X"fc", X"08", 
    X"e6", X"f4", X"fd", X"08", X"e6", X"f4", X"fb", X"08", 
    X"e6", X"f4", X"fe", X"e5", X"0c", X"24", X"0c", X"f8", 
    X"e6", X"52", X"04", X"08", X"e6", X"52", X"05", X"08", 
    X"e6", X"52", X"03", X"08", X"e6", X"52", X"06", X"e5", 
    X"0c", X"24", X"08", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"ec", X"12", X"66", X"a0", 
    X"a3", X"ed", X"12", X"66", X"a0", X"a3", X"eb", X"12", 
    X"66", X"a0", X"a3", X"ee", X"12", X"66", X"a0", X"7f", 
    X"01", X"90", X"00", X"09", X"e0", X"fc", X"a3", X"e0", 
    X"fd", X"a3", X"e0", X"fe", X"74", X"32", X"2c", X"fc", 
    X"e4", X"3d", X"fd", X"8c", X"82", X"8d", X"83", X"8e", 
    X"f0", X"e4", X"12", X"66", X"a0", X"d0", X"e0", X"53", 
    X"e0", X"80", X"e5", X"e0", X"42", X"a8", X"d0", X"e0", 
    X"8f", X"82", X"85", X"0c", X"81", X"d0", X"0c", X"22", 
    X"c0", X"0c", X"e5", X"81", X"f5", X"0c", X"24", X"07", 
    X"f5", X"81", X"af", X"82", X"ae", X"83", X"ad", X"f0", 
    X"e5", X"0c", X"24", X"07", X"f8", X"76", X"01", X"e5", 
    X"0c", X"24", X"04", X"f8", X"a6", X"07", X"08", X"a6", 
    X"06", X"08", X"a6", X"05", X"c0", X"e0", X"c0", X"a8", 
    X"c2", X"af", X"e5", X"0c", X"24", X"f6", X"f8", X"e6", 
    X"08", X"46", X"60", X"52", X"e5", X"0c", X"24", X"f6", 
    X"f8", X"a9", X"0c", X"09", X"e6", X"f7", X"08", X"09", 
    X"e6", X"f7", X"08", X"09", X"e6", X"f7", X"74", X"2e", 
    X"2f", X"fa", X"e4", X"3e", X"fb", X"8d", X"04", X"8a", 
    X"82", X"8b", X"83", X"8c", X"f0", X"12", X"70", X"5a", 
    X"fa", X"a3", X"12", X"70", X"5a", X"fb", X"a3", X"12", 
    X"70", X"5a", X"fc", X"a3", X"12", X"70", X"5a", X"ff", 
    X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"ea", X"12", X"66", X"a0", X"a3", 
    X"eb", X"12", X"66", X"a0", X"a3", X"ec", X"12", X"66", 
    X"a0", X"a3", X"ef", X"12", X"66", X"a0", X"e5", X"0c", 
    X"24", X"04", X"f8", X"74", X"32", X"26", X"fd", X"e4", 
    X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fc", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"74", X"02", 
    X"12", X"66", X"a0", X"e5", X"0c", X"24", X"f9", X"f8", 
    X"e6", X"24", X"fb", X"50", X"03", X"02", X"1b", X"f5", 
    X"e5", X"0c", X"24", X"f9", X"f8", X"e6", X"26", X"26", 
    X"90", X"1a", X"a4", X"73", X"02", X"1b", X"f5", X"02", 
    X"1a", X"b3", X"02", X"1b", X"1f", X"02", X"1b", X"83", 
    X"02", X"1b", X"b6", X"c0", X"04", X"e5", X"0c", X"24", 
    X"04", X"f8", X"a9", X"0c", X"09", X"74", X"2e", X"26", 
    X"f7", X"e4", X"08", X"36", X"09", X"f7", X"08", X"09", 
    X"e6", X"f7", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"fa", X"a3", X"12", X"70", X"5a", X"fb", X"a3", X"12", 
    X"70", X"5a", X"fc", X"a3", X"12", X"70", X"5a", X"ff", 
    X"e5", X"0c", X"24", X"fa", X"f8", X"e6", X"42", X"02", 
    X"08", X"e6", X"42", X"03", X"08", X"e6", X"42", X"04", 
    X"08", X"e6", X"42", X"07", X"a8", X"0c", X"08", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"ea", 
    X"12", X"66", X"a0", X"a3", X"eb", X"12", X"66", X"a0", 
    X"a3", X"ec", X"12", X"66", X"a0", X"a3", X"ef", X"12", 
    X"66", X"a0", X"d0", X"04", X"02", X"1b", X"f5", X"c0", 
    X"04", X"e5", X"0c", X"24", X"04", X"f8", X"a9", X"0c", 
    X"09", X"74", X"2e", X"26", X"f7", X"e4", X"08", X"36", 
    X"09", X"f7", X"08", X"09", X"e6", X"f7", X"a8", X"0c", 
    X"08", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"70", X"5a", X"fa", X"a3", X"12", X"70", 
    X"5a", X"fb", X"a3", X"12", X"70", X"5a", X"fc", X"a3", 
    X"12", X"70", X"5a", X"ff", X"0a", X"ba", X"00", X"09", 
    X"0b", X"bb", X"00", X"05", X"0c", X"bc", X"00", X"01", 
    X"0f", X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"ea", X"12", X"66", X"a0", 
    X"a3", X"eb", X"12", X"66", X"a0", X"a3", X"ec", X"12", 
    X"66", X"a0", X"a3", X"ef", X"12", X"66", X"a0", X"d0", 
    X"04", X"80", X"72", X"e5", X"0c", X"24", X"04", X"f8", 
    X"74", X"2e", X"26", X"fd", X"e4", X"08", X"36", X"fe", 
    X"08", X"86", X"07", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"e5", X"0c", X"24", X"fa", X"f8", X"e6", X"12", 
    X"66", X"a0", X"a3", X"08", X"e6", X"12", X"66", X"a0", 
    X"a3", X"08", X"e6", X"12", X"66", X"a0", X"a3", X"08", 
    X"e6", X"12", X"66", X"a0", X"80", X"3f", X"bc", X"02", 
    X"02", X"80", X"33", X"e5", X"0c", X"24", X"04", X"f8", 
    X"74", X"2e", X"26", X"fd", X"e4", X"08", X"36", X"fe", 
    X"08", X"86", X"07", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"e5", X"0c", X"24", X"fa", X"f8", X"e6", X"12", 
    X"66", X"a0", X"a3", X"08", X"e6", X"12", X"66", X"a0", 
    X"a3", X"08", X"e6", X"12", X"66", X"a0", X"a3", X"08", 
    X"e6", X"12", X"66", X"a0", X"80", X"07", X"e5", X"0c", 
    X"24", X"07", X"f8", X"76", X"00", X"bc", X"01", X"02", 
    X"80", X"03", X"02", X"1c", X"bf", X"e5", X"0c", X"24", 
    X"04", X"f8", X"74", X"03", X"26", X"fd", X"e4", X"08", 
    X"36", X"fe", X"08", X"86", X"07", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"30", X"3b", X"e5", X"0c", 
    X"24", X"04", X"f8", X"74", X"1f", X"26", X"fd", X"e4", 
    X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fc", 
    X"90", X"00", X"69", X"e0", X"c3", X"9c", X"50", X"05", 
    X"90", X"00", X"69", X"ec", X"f0", X"e5", X"0c", X"24", 
    X"04", X"f8", X"a9", X"0c", X"09", X"74", X"03", X"26", 
    X"f7", X"e4", X"08", X"36", X"09", X"f7", X"08", X"09", 
    X"e6", X"f7", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"70", X"5a", X"75", X"f0", X"0c", X"a4", X"24", 
    X"0c", X"fb", X"74", X"00", X"35", X"f0", X"fc", X"7a", 
    X"00", X"c0", X"07", X"c0", X"06", X"c0", X"05", X"a8", 
    X"0c", X"08", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"08", X"e6", X"c0", X"e0", X"8b", X"82", X"8c", 
    X"83", X"8a", X"f0", X"12", X"2c", X"df", X"15", X"81", 
    X"15", X"81", X"15", X"81", X"d0", X"05", X"d0", X"06", 
    X"d0", X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"70", X"5a", X"fd", X"90", X"00", X"09", X"e0", 
    X"fc", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"74", 
    X"1f", X"2c", X"fc", X"e4", X"3e", X"fe", X"8c", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fc", 
    X"c3", X"9d", X"50", X"03", X"12", X"64", X"b5", X"d0", 
    X"e0", X"53", X"e0", X"80", X"e5", X"e0", X"42", X"a8", 
    X"d0", X"e0", X"e5", X"0c", X"24", X"07", X"f8", X"86", 
    X"82", X"85", X"0c", X"81", X"d0", X"0c", X"22", X"c0", 
    X"0c", X"e5", X"81", X"f5", X"0c", X"24", X"07", X"f5", 
    X"81", X"af", X"82", X"ae", X"83", X"ad", X"f0", X"e5", 
    X"0c", X"24", X"07", X"f8", X"76", X"01", X"e5", X"0c", 
    X"24", X"04", X"f8", X"a6", X"07", X"08", X"a6", X"06", 
    X"08", X"a6", X"05", X"e5", X"0c", X"24", X"f6", X"f8", 
    X"e6", X"08", X"46", X"60", X"52", X"e5", X"0c", X"24", 
    X"f6", X"f8", X"a9", X"0c", X"09", X"e6", X"f7", X"08", 
    X"09", X"e6", X"f7", X"08", X"09", X"e6", X"f7", X"74", 
    X"2e", X"2f", X"fa", X"e4", X"3e", X"fb", X"8d", X"04", 
    X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"12", X"70", 
    X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"fb", X"a3", 
    X"12", X"70", X"5a", X"fc", X"a3", X"12", X"70", X"5a", 
    X"ff", X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"ea", X"12", X"66", X"a0", 
    X"a3", X"eb", X"12", X"66", X"a0", X"a3", X"ec", X"12", 
    X"66", X"a0", X"a3", X"ef", X"12", X"66", X"a0", X"e5", 
    X"0c", X"24", X"04", X"f8", X"74", X"32", X"26", X"fd", 
    X"e4", X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"fc", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"74", 
    X"02", X"12", X"66", X"a0", X"e5", X"0c", X"24", X"f9", 
    X"f8", X"e6", X"24", X"fb", X"50", X"03", X"02", X"1e", 
    X"e6", X"e5", X"0c", X"24", X"f9", X"f8", X"e6", X"26", 
    X"26", X"90", X"1d", X"95", X"73", X"02", X"1e", X"e6", 
    X"02", X"1d", X"a4", X"02", X"1e", X"10", X"02", X"1e", 
    X"74", X"02", X"1e", X"a7", X"c0", X"04", X"e5", X"0c", 
    X"24", X"04", X"f8", X"a9", X"0c", X"09", X"74", X"2e", 
    X"26", X"f7", X"e4", X"08", X"36", X"09", X"f7", X"08", 
    X"09", X"e6", X"f7", X"a8", X"0c", X"08", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"70", 
    X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"fb", X"a3", 
    X"12", X"70", X"5a", X"fc", X"a3", X"12", X"70", X"5a", 
    X"ff", X"e5", X"0c", X"24", X"fa", X"f8", X"e6", X"42", 
    X"02", X"08", X"e6", X"42", X"03", X"08", X"e6", X"42", 
    X"04", X"08", X"e6", X"42", X"07", X"a8", X"0c", X"08", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"ea", X"12", X"66", X"a0", X"a3", X"eb", X"12", X"66", 
    X"a0", X"a3", X"ec", X"12", X"66", X"a0", X"a3", X"ef", 
    X"12", X"66", X"a0", X"d0", X"04", X"02", X"1e", X"e6", 
    X"c0", X"04", X"e5", X"0c", X"24", X"04", X"f8", X"a9", 
    X"0c", X"09", X"74", X"2e", X"26", X"f7", X"e4", X"08", 
    X"36", X"09", X"f7", X"08", X"09", X"e6", X"f7", X"a8", 
    X"0c", X"08", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"12", X"70", X"5a", X"fa", X"a3", X"12", 
    X"70", X"5a", X"fb", X"a3", X"12", X"70", X"5a", X"fc", 
    X"a3", X"12", X"70", X"5a", X"ff", X"0a", X"ba", X"00", 
    X"09", X"0b", X"bb", X"00", X"05", X"0c", X"bc", X"00", 
    X"01", X"0f", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"ea", X"12", X"66", 
    X"a0", X"a3", X"eb", X"12", X"66", X"a0", X"a3", X"ec", 
    X"12", X"66", X"a0", X"a3", X"ef", X"12", X"66", X"a0", 
    X"d0", X"04", X"80", X"72", X"e5", X"0c", X"24", X"04", 
    X"f8", X"74", X"2e", X"26", X"fd", X"e4", X"08", X"36", 
    X"fe", X"08", X"86", X"07", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"e5", X"0c", X"24", X"fa", X"f8", X"e6", 
    X"12", X"66", X"a0", X"a3", X"08", X"e6", X"12", X"66", 
    X"a0", X"a3", X"08", X"e6", X"12", X"66", X"a0", X"a3", 
    X"08", X"e6", X"12", X"66", X"a0", X"80", X"3f", X"bc", 
    X"02", X"02", X"80", X"33", X"e5", X"0c", X"24", X"04", 
    X"f8", X"74", X"2e", X"26", X"fd", X"e4", X"08", X"36", 
    X"fe", X"08", X"86", X"07", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"e5", X"0c", X"24", X"fa", X"f8", X"e6", 
    X"12", X"66", X"a0", X"a3", X"08", X"e6", X"12", X"66", 
    X"a0", X"a3", X"08", X"e6", X"12", X"66", X"a0", X"a3", 
    X"08", X"e6", X"12", X"66", X"a0", X"80", X"07", X"e5", 
    X"0c", X"24", X"07", X"f8", X"76", X"00", X"bc", X"01", 
    X"02", X"80", X"03", X"02", X"1f", X"fc", X"90", X"00", 
    X"74", X"e0", X"60", X"03", X"02", X"1f", X"75", X"e5", 
    X"0c", X"24", X"04", X"f8", X"74", X"03", X"26", X"fd", 
    X"e4", X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"30", X"3b", 
    X"e5", X"0c", X"24", X"04", X"f8", X"74", X"1f", X"26", 
    X"fd", X"e4", X"08", X"36", X"fe", X"08", X"86", X"07", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", 
    X"5a", X"fc", X"90", X"00", X"69", X"e0", X"c3", X"9c", 
    X"50", X"05", X"90", X"00", X"69", X"ec", X"f0", X"e5", 
    X"0c", X"24", X"04", X"f8", X"74", X"03", X"26", X"fa", 
    X"e4", X"08", X"36", X"fb", X"08", X"86", X"04", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"75", X"f0", X"0c", X"a4", X"24", X"0c", X"fe", X"74", 
    X"00", X"35", X"f0", X"ff", X"7d", X"00", X"c0", X"02", 
    X"c0", X"03", X"c0", X"04", X"8e", X"82", X"8f", X"83", 
    X"8d", X"f0", X"12", X"2c", X"df", X"15", X"81", X"15", 
    X"81", X"15", X"81", X"80", X"25", X"e5", X"0c", X"24", 
    X"04", X"f8", X"74", X"11", X"26", X"fd", X"e4", X"08", 
    X"36", X"fe", X"08", X"86", X"07", X"c0", X"05", X"c0", 
    X"06", X"c0", X"07", X"90", X"00", X"5a", X"75", X"f0", 
    X"00", X"12", X"2c", X"df", X"15", X"81", X"15", X"81", 
    X"15", X"81", X"e5", X"0c", X"24", X"04", X"f8", X"74", 
    X"1f", X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", 
    X"86", X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"70", X"5a", X"fd", X"90", X"00", X"09", X"e0", 
    X"fc", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"74", 
    X"1f", X"2c", X"fc", X"e4", X"3e", X"fe", X"8c", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fc", 
    X"c3", X"9d", X"50", X"28", X"e5", X"0c", X"24", X"f3", 
    X"f8", X"e6", X"08", X"46", X"60", X"18", X"e5", X"0c", 
    X"24", X"f3", X"f8", X"86", X"05", X"08", X"86", X"06", 
    X"08", X"86", X"07", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"74", X"01", X"12", X"66", X"a0", X"90", X"00", 
    X"6c", X"74", X"01", X"f0", X"e5", X"0c", X"24", X"07", 
    X"f8", X"86", X"82", X"85", X"0c", X"81", X"d0", X"0c", 
    X"22", X"c0", X"0c", X"85", X"81", X"0c", X"c0", X"82", 
    X"c0", X"83", X"c0", X"f0", X"e5", X"81", X"24", X"07", 
    X"f5", X"81", X"a8", X"0c", X"08", X"e5", X"0c", X"24", 
    X"07", X"f9", X"e6", X"f7", X"08", X"09", X"e6", X"f7", 
    X"08", X"09", X"e6", X"f7", X"a8", X"0c", X"08", X"74", 
    X"32", X"26", X"fa", X"e4", X"08", X"36", X"fb", X"08", 
    X"86", X"04", X"8a", X"82", X"8b", X"83", X"8c", X"f0", 
    X"e5", X"0c", X"24", X"0a", X"f8", X"12", X"70", X"5a", 
    X"f6", X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"74", 
    X"02", X"12", X"66", X"a0", X"a8", X"0c", X"08", X"e5", 
    X"0c", X"24", X"04", X"f9", X"74", X"2e", X"26", X"f7", 
    X"e4", X"08", X"36", X"09", X"f7", X"08", X"09", X"e6", 
    X"f7", X"e5", X"0c", X"24", X"04", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"70", 
    X"5a", X"fe", X"a3", X"12", X"70", X"5a", X"fd", X"a3", 
    X"12", X"70", X"5a", X"fc", X"a3", X"12", X"70", X"5a", 
    X"ff", X"0e", X"be", X"00", X"09", X"0d", X"bd", X"00", 
    X"05", X"0c", X"bc", X"00", X"01", X"0f", X"e5", X"0c", 
    X"24", X"04", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"ee", X"12", X"66", X"a0", X"a3", 
    X"ed", X"12", X"66", X"a0", X"a3", X"ec", X"12", X"66", 
    X"a0", X"a3", X"ef", X"12", X"66", X"a0", X"e5", X"0c", 
    X"24", X"0a", X"f8", X"b6", X"01", X"02", X"80", X"03", 
    X"02", X"21", X"db", X"90", X"00", X"74", X"e0", X"60", 
    X"03", X"02", X"21", X"56", X"a8", X"0c", X"08", X"74", 
    X"03", X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", 
    X"86", X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"30", X"3b", X"a8", X"0c", X"08", X"74", X"1f", 
    X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", X"86", 
    X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"70", X"5a", X"ff", X"90", X"00", X"69", X"e0", X"c3", 
    X"9f", X"50", X"05", X"90", X"00", X"69", X"ef", X"f0", 
    X"e5", X"0c", X"24", X"07", X"f8", X"74", X"03", X"26", 
    X"fd", X"e4", X"08", X"36", X"fe", X"08", X"86", X"07", 
    X"e5", X"0c", X"24", X"07", X"f8", X"74", X"1f", X"26", 
    X"fa", X"e4", X"08", X"36", X"fb", X"08", X"86", X"04", 
    X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"12", X"70", 
    X"5a", X"75", X"f0", X"0c", X"a4", X"24", X"0c", X"fb", 
    X"74", X"00", X"35", X"f0", X"fc", X"7a", X"00", X"c0", 
    X"05", X"c0", X"06", X"c0", X"07", X"8b", X"82", X"8c", 
    X"83", X"8a", X"f0", X"12", X"2c", X"df", X"15", X"81", 
    X"15", X"81", X"15", X"81", X"80", X"23", X"a8", X"0c", 
    X"08", X"74", X"11", X"26", X"fd", X"e4", X"08", X"36", 
    X"fe", X"08", X"86", X"07", X"c0", X"05", X"c0", X"06", 
    X"c0", X"07", X"90", X"00", X"5a", X"75", X"f0", X"00", 
    X"12", X"2c", X"df", X"15", X"81", X"15", X"81", X"15", 
    X"81", X"e5", X"0c", X"24", X"07", X"f8", X"74", X"1f", 
    X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", X"86", 
    X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"70", X"5a", X"fd", X"90", X"00", X"09", X"e0", X"fc", 
    X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"74", X"1f", 
    X"2c", X"fc", X"e4", X"3e", X"fe", X"8c", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fc", X"c3", 
    X"9d", X"50", X"28", X"e5", X"0c", X"24", X"fb", X"f8", 
    X"e6", X"08", X"46", X"60", X"18", X"e5", X"0c", X"24", 
    X"fb", X"f8", X"86", X"05", X"08", X"86", X"06", X"08", 
    X"86", X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"74", X"01", X"12", X"66", X"a0", X"90", X"00", X"6c", 
    X"74", X"01", X"f0", X"85", X"0c", X"81", X"d0", X"0c", 
    X"22", X"ad", X"82", X"ae", X"83", X"af", X"f0", X"ed", 
    X"4e", X"70", X"0d", X"90", X"00", X"09", X"e0", X"fa", 
    X"a3", X"e0", X"fb", X"a3", X"e0", X"fc", X"80", X"06", 
    X"8d", X"02", X"8e", X"03", X"8f", X"04", X"c0", X"e0", 
    X"c0", X"a8", X"c2", X"af", X"74", X"32", X"2a", X"fd", 
    X"e4", X"3b", X"fe", X"8c", X"07", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fc", X"bc", 
    X"02", X"0e", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"e4", X"12", X"66", X"a0", X"7f", X"01", X"80", X"02", 
    X"7f", X"00", X"d0", X"e0", X"53", X"e0", X"80", X"e5", 
    X"e0", X"42", X"a8", X"d0", X"e0", X"8f", X"82", X"22", 
    X"c0", X"0c", X"85", X"81", X"0c", X"c0", X"82", X"c0", 
    X"83", X"e5", X"81", X"24", X"04", X"f5", X"81", X"90", 
    X"00", X"67", X"e0", X"fc", X"a3", X"e0", X"fd", X"e5", 
    X"0c", X"24", X"05", X"f8", X"a6", X"04", X"08", X"a6", 
    X"05", X"90", X"00", X"09", X"e0", X"fa", X"a3", X"e0", 
    X"fb", X"a3", X"e0", X"ff", X"74", X"03", X"2a", X"fa", 
    X"e4", X"3b", X"fb", X"8a", X"82", X"8b", X"83", X"8f", 
    X"f0", X"12", X"30", X"3b", X"e5", X"0c", X"24", X"05", 
    X"f8", X"a9", X"0c", X"09", X"e7", X"26", X"fe", X"09", 
    X"e7", X"08", X"36", X"ff", X"e5", X"0c", X"24", X"03", 
    X"f8", X"a6", X"06", X"08", X"a6", X"07", X"90", X"00", 
    X"09", X"e0", X"fa", X"a3", X"e0", X"fb", X"a3", X"e0", 
    X"fd", X"74", X"03", X"2a", X"fa", X"e4", X"3b", X"fb", 
    X"8a", X"82", X"8b", X"83", X"8d", X"f0", X"e5", X"0c", 
    X"24", X"03", X"f8", X"e6", X"12", X"66", X"a0", X"a3", 
    X"08", X"e6", X"12", X"66", X"a0", X"e5", X"0c", X"24", 
    X"03", X"f8", X"e5", X"0c", X"24", X"05", X"f9", X"c3", 
    X"e6", X"97", X"08", X"e6", X"09", X"97", X"50", X"36", 
    X"90", X"00", X"09", X"e0", X"fb", X"a3", X"e0", X"fc", 
    X"a3", X"e0", X"fd", X"74", X"03", X"2b", X"fb", X"e4", 
    X"3c", X"fe", X"8d", X"07", X"90", X"00", X"57", X"e0", 
    X"fa", X"a3", X"e0", X"fc", X"a3", X"e0", X"fd", X"c0", 
    X"03", X"c0", X"06", X"c0", X"07", X"8a", X"82", X"8c", 
    X"83", X"8d", X"f0", X"12", X"2e", X"3d", X"15", X"81", 
    X"15", X"81", X"15", X"81", X"80", X"55", X"90", X"00", 
    X"09", X"e0", X"fb", X"a3", X"e0", X"fc", X"a3", X"e0", 
    X"fd", X"74", X"03", X"2b", X"fb", X"e4", X"3c", X"fc", 
    X"90", X"00", X"54", X"e0", X"fa", X"a3", X"e0", X"fe", 
    X"a3", X"e0", X"ff", X"c0", X"03", X"c0", X"04", X"c0", 
    X"05", X"8a", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"2e", X"3d", X"15", X"81", X"15", X"81", X"15", X"81", 
    X"90", X"00", X"6f", X"e0", X"fe", X"a3", X"e0", X"ff", 
    X"e5", X"0c", X"24", X"03", X"f8", X"c3", X"e6", X"9e", 
    X"08", X"e6", X"9f", X"50", X"0e", X"e5", X"0c", X"24", 
    X"03", X"f8", X"90", X"00", X"6f", X"e6", X"f0", X"08", 
    X"e6", X"a3", X"f0", X"85", X"0c", X"81", X"d0", X"0c", 
    X"22", X"90", X"00", X"0e", X"12", X"61", X"84", X"ad", 
    X"82", X"ae", X"83", X"af", X"f0", X"ed", X"4e", X"60", 
    X"2c", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"e4", 
    X"12", X"66", X"a0", X"a3", X"12", X"66", X"a0", X"74", 
    X"02", X"2d", X"fa", X"e4", X"3e", X"fb", X"8f", X"04", 
    X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"c0", X"07", 
    X"c0", X"06", X"c0", X"05", X"12", X"2b", X"dd", X"d0", 
    X"05", X"d0", X"06", X"d0", X"07", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"22", X"c0", X"0c", X"85", X"81", 
    X"0c", X"c0", X"82", X"c0", X"83", X"c0", X"f0", X"e5", 
    X"81", X"24", X"05", X"f5", X"81", X"a8", X"0c", X"08", 
    X"e5", X"0c", X"24", X"04", X"f9", X"e6", X"f7", X"08", 
    X"09", X"e6", X"f7", X"08", X"09", X"e6", X"f7", X"12", 
    X"09", X"4a", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"ff", X"a3", X"12", X"70", X"5a", X"fe", X"c0", X"07", 
    X"c0", X"06", X"e5", X"0c", X"24", X"fc", X"f8", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"a8", X"0c", 
    X"08", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"28", X"28", X"15", X"81", X"15", X"81", 
    X"d0", X"06", X"d0", X"07", X"e5", X"0c", X"24", X"fc", 
    X"f8", X"e6", X"4f", X"fa", X"08", X"e6", X"4e", X"fc", 
    X"e5", X"0c", X"24", X"fa", X"f8", X"e6", X"52", X"02", 
    X"08", X"e6", X"52", X"04", X"e5", X"0c", X"24", X"fa", 
    X"f8", X"e6", X"b5", X"02", X"07", X"08", X"e6", X"b5", 
    X"04", X"02", X"80", X"02", X"80", X"51", X"e5", X"0c", 
    X"24", X"fc", X"f8", X"e6", X"4f", X"fb", X"08", X"e6", 
    X"4e", X"fc", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"fa", X"a3", X"12", X"70", X"5a", X"ff", X"e5", X"0c", 
    X"24", X"fa", X"f8", X"e6", X"f4", X"fd", X"08", X"e6", 
    X"f4", X"fe", X"ed", X"52", X"02", X"ee", X"52", X"07", 
    X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"ea", X"12", X"66", X"a0", X"a3", 
    X"ef", X"12", X"66", X"a0", X"e5", X"0c", X"24", X"f8", 
    X"f8", X"e4", X"f6", X"08", X"f6", X"80", X"5d", X"e5", 
    X"0c", X"24", X"f8", X"f8", X"e6", X"08", X"46", X"60", 
    X"3f", X"e5", X"0c", X"24", X"fa", X"f8", X"86", X"06", 
    X"74", X"05", X"08", X"46", X"fc", X"a8", X"0c", X"08", 
    X"74", X"02", X"26", X"fa", X"e4", X"08", X"36", X"fd", 
    X"08", X"86", X"07", X"e5", X"0c", X"24", X"f8", X"f8", 
    X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"c0", 
    X"06", X"c0", X"04", X"8a", X"82", X"8d", X"83", X"8f", 
    X"f0", X"12", X"0f", X"da", X"e5", X"81", X"24", X"fc", 
    X"f5", X"81", X"7b", X"00", X"7c", X"00", X"80", X"14", 
    X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"70", X"5a", X"fb", X"a3", 
    X"12", X"70", X"5a", X"fc", X"c0", X"04", X"c0", X"03", 
    X"12", X"09", X"52", X"af", X"82", X"d0", X"03", X"d0", 
    X"04", X"e5", X"0c", X"24", X"f8", X"f8", X"e6", X"08", 
    X"46", X"70", X"03", X"02", X"25", X"98", X"ef", X"70", 
    X"03", X"12", X"64", X"b5", X"12", X"15", X"59", X"ae", 
    X"82", X"af", X"83", X"e5", X"0c", X"24", X"07", X"f8", 
    X"a6", X"06", X"08", X"a6", X"07", X"e5", X"0c", X"24", 
    X"07", X"f8", X"08", X"e6", X"30", X"e1", X"03", X"02", 
    X"25", X"8f", X"c0", X"e0", X"c0", X"a8", X"c2", X"af", 
    X"e5", X"0c", X"24", X"04", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"fa", X"a3", X"12", X"70", X"5a", X"fd", X"e5", X"0c", 
    X"24", X"07", X"f8", X"a6", X"02", X"08", X"a6", X"05", 
    X"e5", X"0c", X"24", X"07", X"f8", X"e5", X"0c", X"24", 
    X"fa", X"f9", X"e7", X"56", X"fe", X"09", X"e7", X"08", 
    X"56", X"ff", X"e5", X"0c", X"24", X"fa", X"f8", X"e6", 
    X"b5", X"06", X"07", X"08", X"e6", X"b5", X"07", X"02", 
    X"80", X"02", X"80", X"28", X"e5", X"0c", X"24", X"fa", 
    X"f8", X"e6", X"f4", X"fe", X"08", X"e6", X"f4", X"ff", 
    X"ee", X"52", X"02", X"ef", X"52", X"05", X"e5", X"0c", 
    X"24", X"04", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"ea", X"12", X"66", X"a0", X"a3", 
    X"ed", X"12", X"66", X"a0", X"d0", X"e0", X"53", X"e0", 
    X"80", X"e5", X"e0", X"42", X"a8", X"d0", X"e0", X"e5", 
    X"0c", X"24", X"07", X"f8", X"86", X"03", X"7c", X"00", 
    X"8b", X"82", X"8c", X"83", X"85", X"0c", X"81", X"d0", 
    X"0c", X"22", X"c0", X"0c", X"85", X"81", X"0c", X"c0", 
    X"82", X"c0", X"83", X"c0", X"f0", X"05", X"81", X"05", 
    X"81", X"05", X"81", X"a8", X"0c", X"08", X"e5", X"0c", 
    X"24", X"04", X"f9", X"e6", X"f7", X"08", X"09", X"e6", 
    X"f7", X"08", X"09", X"e6", X"f7", X"7f", X"00", X"7e", 
    X"00", X"c0", X"07", X"c0", X"06", X"12", X"09", X"4a", 
    X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"70", X"5a", X"fd", X"a3", 
    X"12", X"70", X"5a", X"fa", X"c0", X"05", X"c0", X"02", 
    X"e5", X"0c", X"24", X"fa", X"f8", X"e6", X"c0", X"e0", 
    X"e5", X"0c", X"24", X"fc", X"f8", X"e6", X"c0", X"e0", 
    X"08", X"e6", X"c0", X"e0", X"8d", X"82", X"8a", X"83", 
    X"12", X"2b", X"92", X"ac", X"82", X"15", X"81", X"15", 
    X"81", X"15", X"81", X"d0", X"02", X"d0", X"05", X"d0", 
    X"06", X"d0", X"07", X"ec", X"60", X"5c", X"8d", X"03", 
    X"8a", X"04", X"e5", X"0c", X"24", X"f8", X"f8", X"e4", 
    X"f6", X"08", X"f6", X"e5", X"0c", X"24", X"fb", X"f8", 
    X"e6", X"70", X"03", X"02", X"26", X"d8", X"c0", X"03", 
    X"c0", X"04", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"fa", X"a3", X"12", X"70", X"5a", X"fc", X"e5", X"0c", 
    X"24", X"fc", X"f8", X"e6", X"f4", X"fb", X"08", X"e6", 
    X"f4", X"ff", X"eb", X"52", X"02", X"ef", X"52", X"04", 
    X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"ea", X"12", X"66", X"a0", X"a3", 
    X"ec", X"12", X"66", X"a0", X"d0", X"04", X"d0", X"03", 
    X"80", X"66", X"e5", X"0c", X"24", X"f8", X"f8", X"e6", 
    X"08", X"46", X"70", X"06", X"8d", X"03", X"8a", X"04", 
    X"80", X"56", X"e5", X"0c", X"24", X"fb", X"f8", X"e6", 
    X"60", X"04", X"7f", X"00", X"7e", X"01", X"e5", X"0c", 
    X"24", X"fa", X"f8", X"e6", X"60", X"03", X"43", X"06", 
    X"04", X"e5", X"0c", X"24", X"fc", X"f8", X"ef", X"46", 
    X"fc", X"ee", X"08", X"46", X"fe", X"e5", X"0c", X"24", 
    X"04", X"f8", X"74", X"02", X"26", X"fa", X"e4", X"08", 
    X"36", X"fd", X"08", X"86", X"07", X"e5", X"0c", X"24", 
    X"f8", X"f8", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"c0", X"04", X"c0", X"06", X"8a", X"82", X"8d", 
    X"83", X"8f", X"f0", X"12", X"0f", X"da", X"e5", X"81", 
    X"24", X"fc", X"f5", X"81", X"7b", X"00", X"7c", X"00", 
    X"c0", X"04", X"c0", X"03", X"12", X"09", X"52", X"af", 
    X"82", X"d0", X"03", X"d0", X"04", X"e5", X"0c", X"24", 
    X"f8", X"f8", X"e6", X"08", X"46", X"70", X"03", X"02", 
    X"27", X"ad", X"ef", X"70", X"03", X"12", X"64", X"b5", 
    X"12", X"15", X"59", X"ae", X"82", X"e5", X"83", X"ff", 
    X"30", X"e1", X"03", X"02", X"27", X"a9", X"c0", X"e0", 
    X"c0", X"a8", X"c2", X"af", X"e5", X"0c", X"24", X"04", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"70", X"5a", X"fe", X"a3", X"12", X"70", 
    X"5a", X"ff", X"c0", X"07", X"c0", X"06", X"e5", X"0c", 
    X"24", X"fa", X"f8", X"e6", X"c0", X"e0", X"e5", X"0c", 
    X"24", X"fc", X"f8", X"e6", X"c0", X"e0", X"08", X"e6", 
    X"c0", X"e0", X"8e", X"82", X"8f", X"83", X"12", X"2b", 
    X"92", X"ad", X"82", X"15", X"81", X"15", X"81", X"15", 
    X"81", X"d0", X"06", X"d0", X"07", X"ed", X"60", X"4e", 
    X"e5", X"0c", X"24", X"fb", X"f8", X"e6", X"60", X"46", 
    X"c0", X"06", X"c0", X"07", X"e5", X"0c", X"24", X"04", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"70", X"5a", X"fa", X"a3", X"12", X"70", 
    X"5a", X"fd", X"e5", X"0c", X"24", X"fc", X"f8", X"e6", 
    X"f4", X"fe", X"08", X"e6", X"f4", X"ff", X"ee", X"52", 
    X"02", X"ef", X"52", X"05", X"e5", X"0c", X"24", X"04", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"ea", X"12", X"66", X"a0", X"a3", X"ed", X"12", 
    X"66", X"a0", X"d0", X"07", X"d0", X"06", X"d0", X"e0", 
    X"53", X"e0", X"80", X"e5", X"e0", X"42", X"a8", X"d0", 
    X"e0", X"8e", X"03", X"7c", X"00", X"8b", X"82", X"8c", 
    X"83", X"85", X"0c", X"81", X"d0", X"0c", X"22", X"c0", 
    X"0c", X"85", X"81", X"0c", X"c0", X"82", X"c0", X"83", 
    X"c0", X"f0", X"c0", X"e0", X"c0", X"a8", X"c2", X"af", 
    X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"70", X"5a", X"fe", X"a3", 
    X"12", X"70", X"5a", X"fd", X"8e", X"02", X"8d", X"04", 
    X"e5", X"0c", X"24", X"fc", X"f8", X"e6", X"f4", X"fb", 
    X"08", X"e6", X"f4", X"ff", X"ee", X"52", X"03", X"ed", 
    X"52", X"07", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"eb", X"12", X"66", 
    X"a0", X"a3", X"ef", X"12", X"66", X"a0", X"d0", X"e0", 
    X"53", X"e0", X"80", X"e5", X"e0", X"42", X"a8", X"d0", 
    X"e0", X"8a", X"82", X"8c", X"83", X"85", X"0c", X"81", 
    X"d0", X"0c", X"22", X"12", X"70", X"5a", X"fd", X"a3", 
    X"12", X"70", X"5a", X"8d", X"82", X"f5", X"83", X"22", 
    X"c0", X"0c", X"e5", X"81", X"f5", X"0c", X"24", X"10", 
    X"f5", X"81", X"aa", X"82", X"ab", X"83", X"ac", X"f0", 
    X"e5", X"0c", X"24", X"0a", X"f8", X"e4", X"f6", X"08", 
    X"f6", X"e5", X"0c", X"24", X"0e", X"f8", X"a6", X"02", 
    X"08", X"a6", X"03", X"08", X"a6", X"04", X"e5", X"0c", 
    X"24", X"07", X"f8", X"74", X"02", X"2a", X"f6", X"e4", 
    X"3b", X"08", X"f6", X"08", X"a6", X"04", X"e5", X"0c", 
    X"24", X"07", X"f8", X"74", X"04", X"26", X"fd", X"e4", 
    X"08", X"36", X"fe", X"08", X"86", X"07", X"e5", X"0c", 
    X"24", X"04", X"f8", X"a6", X"05", X"08", X"a6", X"06", 
    X"08", X"a6", X"07", X"c0", X"04", X"c0", X"03", X"c0", 
    X"02", X"12", X"09", X"4a", X"d0", X"02", X"d0", X"03", 
    X"d0", X"04", X"e5", X"0c", X"24", X"07", X"f8", X"74", 
    X"06", X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", 
    X"86", X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"a8", X"0c", X"08", X"12", X"70", X"5a", X"f6", X"a3", 
    X"12", X"70", X"5a", X"08", X"f6", X"a3", X"12", X"70", 
    X"5a", X"08", X"f6", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"12", X"70", X"5a", X"fe", X"a3", X"12", X"70", 
    X"5a", X"ff", X"e5", X"0c", X"24", X"fc", X"f8", X"e6", 
    X"42", X"06", X"08", X"e6", X"42", X"07", X"8a", X"82", 
    X"8b", X"83", X"8c", X"f0", X"ee", X"12", X"66", X"a0", 
    X"a3", X"ef", X"12", X"66", X"a0", X"a8", X"0c", X"08", 
    X"e5", X"0c", X"24", X"04", X"f9", X"e7", X"c0", X"e0", 
    X"09", X"e7", X"c0", X"e0", X"09", X"e7", X"c0", X"e0", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"12", X"00", X"11", X"15", X"81", X"15", X"81", X"15", 
    X"81", X"70", X"03", X"02", X"2a", X"2e", X"a8", X"0c", 
    X"08", X"74", X"02", X"26", X"fd", X"e4", X"08", X"36", 
    X"fe", X"08", X"86", X"07", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"70", X"5a", X"fd", X"a3", X"12", 
    X"70", X"5a", X"fe", X"a3", X"12", X"70", X"5a", X"ff", 
    X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"70", X"5a", X"fb", X"a3", 
    X"12", X"70", X"5a", X"fc", X"7a", X"00", X"e5", X"0c", 
    X"24", X"0c", X"f8", X"76", X"00", X"08", X"a6", X"04", 
    X"7c", X"00", X"e5", X"0c", X"24", X"0c", X"f8", X"08", 
    X"e6", X"20", X"e2", X"30", X"c0", X"05", X"c0", X"06", 
    X"c0", X"07", X"e5", X"0c", X"24", X"0e", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"12", 
    X"70", X"5a", X"fe", X"a3", X"12", X"70", X"5a", X"ff", 
    X"eb", X"52", X"06", X"ec", X"52", X"07", X"ee", X"4f", 
    X"d0", X"07", X"d0", X"06", X"d0", X"05", X"60", X"40", 
    X"7a", X"01", X"80", X"3c", X"c0", X"05", X"c0", X"06", 
    X"c0", X"07", X"e5", X"0c", X"24", X"0e", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"12", 
    X"70", X"5a", X"fe", X"a3", X"12", X"70", X"5a", X"ff", 
    X"eb", X"52", X"06", X"ec", X"52", X"07", X"ee", X"b5", 
    X"03", X"06", X"ef", X"b5", X"04", X"02", X"80", X"08", 
    X"d0", X"07", X"d0", X"06", X"d0", X"05", X"80", X"08", 
    X"d0", X"07", X"d0", X"06", X"d0", X"05", X"7a", X"01", 
    X"ea", X"60", X"5d", X"e5", X"0c", X"24", X"0c", X"f8", 
    X"08", X"e6", X"30", X"e0", X"0c", X"e5", X"0c", X"24", 
    X"0a", X"f8", X"eb", X"46", X"f6", X"ec", X"08", X"46", 
    X"f6", X"c0", X"05", X"c0", X"06", X"c0", X"07", X"e5", 
    X"0c", X"24", X"0e", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", X"fe", 
    X"a3", X"12", X"70", X"5a", X"ff", X"43", X"07", X"02", 
    X"c0", X"07", X"c0", X"06", X"c0", X"05", X"c0", X"06", 
    X"c0", X"07", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"11", X"b5", 
    X"15", X"81", X"15", X"81", X"d0", X"05", X"d0", X"06", 
    X"d0", X"07", X"d0", X"07", X"d0", X"06", X"d0", X"05", 
    X"a8", X"0c", X"08", X"a6", X"05", X"08", X"a6", X"06", 
    X"08", X"a6", X"07", X"02", X"28", X"dd", X"e5", X"0c", 
    X"24", X"0e", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"70", X"5a", X"fe", X"a3", 
    X"12", X"70", X"5a", X"ff", X"e5", X"0c", X"24", X"0a", 
    X"f8", X"e6", X"f4", X"fc", X"08", X"e6", X"f4", X"fd", 
    X"ec", X"52", X"06", X"ed", X"52", X"07", X"e5", X"0c", 
    X"24", X"0e", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"ee", X"12", X"66", X"a0", X"a3", 
    X"ef", X"12", X"66", X"a0", X"12", X"09", X"52", X"e5", 
    X"0c", X"24", X"0e", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", X"fe", 
    X"a3", X"12", X"70", X"5a", X"ff", X"8e", X"82", X"8f", 
    X"83", X"85", X"0c", X"81", X"d0", X"0c", X"22", X"c0", 
    X"0c", X"85", X"81", X"0c", X"05", X"81", X"05", X"81", 
    X"05", X"81", X"ad", X"82", X"ae", X"83", X"af", X"f0", 
    X"a8", X"0c", X"08", X"a6", X"05", X"08", X"a6", X"06", 
    X"08", X"a6", X"07", X"74", X"02", X"2d", X"fd", X"e4", 
    X"3e", X"fe", X"c0", X"07", X"c0", X"06", X"c0", X"05", 
    X"12", X"09", X"4a", X"d0", X"05", X"d0", X"06", X"d0", 
    X"07", X"74", X"06", X"2d", X"fa", X"e4", X"3e", X"fb", 
    X"8f", X"04", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"70", X"5a", X"60", X"4e", X"c0", X"05", X"c0", 
    X"06", X"c0", X"07", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"12", X"70", X"5a", X"fd", X"a3", X"12", X"70", 
    X"5a", X"fe", X"a3", X"12", X"70", X"5a", X"ff", X"c0", 
    X"07", X"c0", X"06", X"c0", X"05", X"c0", X"04", X"c0", 
    X"03", X"c0", X"02", X"e4", X"c0", X"e0", X"74", X"02", 
    X"c0", X"e0", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"11", X"b5", X"15", X"81", X"15", X"81", X"d0", 
    X"02", X"d0", X"03", X"d0", X"04", X"d0", X"05", X"d0", 
    X"06", X"d0", X"07", X"d0", X"07", X"d0", X"06", X"d0", 
    X"05", X"80", X"a7", X"a8", X"0c", X"08", X"86", X"02", 
    X"08", X"86", X"03", X"08", X"86", X"04", X"8a", X"82", 
    X"8b", X"83", X"8c", X"f0", X"12", X"62", X"2d", X"12", 
    X"09", X"52", X"85", X"0c", X"81", X"d0", X"0c", X"22", 
    X"c0", X"0c", X"85", X"81", X"0c", X"ad", X"82", X"ae", 
    X"83", X"af", X"f0", X"e5", X"0c", X"24", X"fa", X"f8", 
    X"86", X"03", X"08", X"86", X"04", X"c0", X"03", X"c0", 
    X"04", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"28", X"28", X"15", X"81", X"15", X"81", X"d0", X"0c", 
    X"22", X"c0", X"0c", X"85", X"81", X"0c", X"ad", X"82", 
    X"ae", X"83", X"af", X"f0", X"e5", X"0c", X"24", X"fa", 
    X"f8", X"86", X"03", X"08", X"86", X"04", X"c0", X"03", 
    X"c0", X"04", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"27", X"b7", X"15", X"81", X"15", X"81", X"d0", 
    X"0c", X"22", X"c0", X"0c", X"85", X"81", X"0c", X"ae", 
    X"82", X"af", X"83", X"7d", X"00", X"e5", X"0c", X"24", 
    X"fb", X"f8", X"e6", X"70", X"13", X"e5", X"0c", X"24", 
    X"fc", X"f8", X"e6", X"5e", X"fb", X"08", X"e6", X"5f", 
    X"fc", X"4b", X"60", X"24", X"7d", X"01", X"80", X"20", 
    X"e5", X"0c", X"24", X"fc", X"f8", X"e6", X"52", X"06", 
    X"08", X"e6", X"52", X"07", X"e5", X"0c", X"24", X"fc", 
    X"f8", X"e6", X"b5", X"06", X"07", X"08", X"e6", X"b5", 
    X"07", X"02", X"80", X"02", X"80", X"02", X"7d", X"01", 
    X"8d", X"82", X"d0", X"0c", X"22", X"c0", X"0c", X"85", 
    X"81", X"0c", X"c0", X"82", X"c0", X"83", X"c0", X"f0", 
    X"05", X"81", X"05", X"81", X"05", X"81", X"a8", X"0c", 
    X"08", X"74", X"01", X"26", X"ff", X"e4", X"08", X"36", 
    X"fb", X"08", X"86", X"02", X"a8", X"0c", X"08", X"e5", 
    X"0c", X"24", X"04", X"f9", X"74", X"04", X"26", X"f7", 
    X"e4", X"08", X"36", X"09", X"f7", X"08", X"09", X"e6", 
    X"f7", X"e5", X"0c", X"24", X"04", X"f8", X"86", X"04", 
    X"08", X"86", X"05", X"08", X"86", X"06", X"8f", X"82", 
    X"8b", X"83", X"8a", X"f0", X"ec", X"12", X"66", X"a0", 
    X"a3", X"ed", X"12", X"66", X"a0", X"a3", X"ee", X"12", 
    X"66", X"a0", X"e5", X"0c", X"24", X"04", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"74", 
    X"ff", X"12", X"66", X"a0", X"a3", X"12", X"66", X"a0", 
    X"e5", X"0c", X"24", X"04", X"f8", X"74", X"02", X"26", 
    X"ff", X"e4", X"08", X"36", X"fd", X"08", X"86", X"04", 
    X"e5", X"0c", X"24", X"04", X"f8", X"86", X"02", X"08", 
    X"86", X"03", X"08", X"86", X"06", X"8f", X"82", X"8d", 
    X"83", X"8c", X"f0", X"ea", X"12", X"66", X"a0", X"a3", 
    X"eb", X"12", X"66", X"a0", X"a3", X"ee", X"12", X"66", 
    X"a0", X"e5", X"0c", X"24", X"04", X"f8", X"74", X"05", 
    X"26", X"ff", X"e4", X"08", X"36", X"fd", X"08", X"86", 
    X"04", X"e5", X"0c", X"24", X"04", X"f8", X"86", X"02", 
    X"08", X"86", X"03", X"08", X"86", X"06", X"8f", X"82", 
    X"8d", X"83", X"8c", X"f0", X"ea", X"12", X"66", X"a0", 
    X"a3", X"eb", X"12", X"66", X"a0", X"a3", X"ee", X"12", 
    X"66", X"a0", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"e4", X"12", X"66", 
    X"a0", X"85", X"0c", X"81", X"d0", X"0c", X"22", X"ad", 
    X"82", X"ae", X"83", X"af", X"f0", X"74", X"0b", X"2d", 
    X"fd", X"e4", X"3e", X"fe", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"e4", X"12", X"66", X"a0", X"a3", X"12", 
    X"66", X"a0", X"a3", X"12", X"66", X"a0", X"22", X"c0", 
    X"0c", X"85", X"81", X"0c", X"c0", X"82", X"c0", X"83", 
    X"c0", X"f0", X"e5", X"81", X"24", X"09", X"f5", X"81", 
    X"a8", X"0c", X"08", X"74", X"01", X"26", X"fa", X"e4", 
    X"08", X"36", X"fb", X"08", X"86", X"04", X"8a", X"82", 
    X"8b", X"83", X"8c", X"f0", X"e5", X"0c", X"24", X"0a", 
    X"f8", X"12", X"70", X"5a", X"f6", X"a3", X"12", X"70", 
    X"5a", X"08", X"f6", X"a3", X"12", X"70", X"5a", X"08", 
    X"f6", X"e5", X"0c", X"24", X"fb", X"f8", X"86", X"02", 
    X"08", X"86", X"03", X"08", X"86", X"04", X"74", X"02", 
    X"2a", X"fd", X"e4", X"3b", X"fe", X"8c", X"07", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"e5", X"0c", X"24", 
    X"0a", X"f8", X"e6", X"12", X"66", X"a0", X"a3", X"08", 
    X"e6", X"12", X"66", X"a0", X"a3", X"08", X"e6", X"12", 
    X"66", X"a0", X"e5", X"0c", X"24", X"04", X"f8", X"74", 
    X"05", X"2a", X"f6", X"e4", X"3b", X"08", X"f6", X"08", 
    X"a6", X"04", X"e5", X"0c", X"24", X"0a", X"f8", X"e5", 
    X"0c", X"24", X"07", X"f9", X"74", X"05", X"26", X"f7", 
    X"e4", X"08", X"36", X"09", X"f7", X"08", X"09", X"e6", 
    X"f7", X"e5", X"0c", X"24", X"07", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"70", 
    X"5a", X"fd", X"a3", X"12", X"70", X"5a", X"fe", X"a3", 
    X"12", X"70", X"5a", X"ff", X"e5", X"0c", X"24", X"04", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"ed", X"12", X"66", X"a0", X"a3", X"ee", X"12", 
    X"66", X"a0", X"a3", X"ef", X"12", X"66", X"a0", X"e5", 
    X"0c", X"24", X"07", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", X"fd", 
    X"a3", X"12", X"70", X"5a", X"fe", X"a3", X"12", X"70", 
    X"5a", X"ff", X"74", X"02", X"2d", X"fd", X"e4", X"3e", 
    X"fe", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"ea", 
    X"12", X"66", X"a0", X"a3", X"eb", X"12", X"66", X"a0", 
    X"a3", X"ec", X"12", X"66", X"a0", X"e5", X"0c", X"24", 
    X"07", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"ea", X"12", X"66", X"a0", X"a3", X"eb", 
    X"12", X"66", X"a0", X"a3", X"ec", X"12", X"66", X"a0", 
    X"74", X"0b", X"2a", X"fa", X"e4", X"3b", X"fb", X"8a", 
    X"82", X"8b", X"83", X"8c", X"f0", X"a8", X"0c", X"08", 
    X"e6", X"12", X"66", X"a0", X"a3", X"08", X"e6", X"12", 
    X"66", X"a0", X"a3", X"08", X"e6", X"12", X"66", X"a0", 
    X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"70", X"5a", X"ff", X"0f", 
    X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"ef", X"12", X"66", X"a0", X"85", 
    X"0c", X"81", X"d0", X"0c", X"22", X"c0", X"0c", X"85", 
    X"81", X"0c", X"c0", X"82", X"c0", X"83", X"c0", X"f0", 
    X"e5", X"81", X"24", X"0b", X"f5", X"81", X"e5", X"0c", 
    X"24", X"fb", X"f8", X"86", X"02", X"08", X"86", X"03", 
    X"08", X"86", X"04", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"e5", X"0c", X"24", X"0d", X"f8", X"12", X"70", 
    X"5a", X"f6", X"a3", X"12", X"70", X"5a", X"08", X"f6", 
    X"e5", X"0c", X"24", X"0d", X"f8", X"b6", X"ff", X"43", 
    X"08", X"b6", X"ff", X"3f", X"c0", X"02", X"c0", X"03", 
    X"c0", X"04", X"a8", X"0c", X"08", X"74", X"04", X"26", 
    X"fa", X"e4", X"08", X"36", X"fb", X"08", X"86", X"04", 
    X"74", X"05", X"2a", X"fa", X"e4", X"3b", X"fb", X"8a", 
    X"82", X"8b", X"83", X"8c", X"f0", X"e5", X"0c", X"24", 
    X"0a", X"f8", X"12", X"70", X"5a", X"f6", X"a3", X"12", 
    X"70", X"5a", X"08", X"f6", X"a3", X"12", X"70", X"5a", 
    X"08", X"f6", X"d0", X"04", X"d0", X"03", X"d0", X"02", 
    X"02", X"2f", X"3f", X"a8", X"0c", X"08", X"74", X"04", 
    X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", X"86", 
    X"07", X"e5", X"0c", X"24", X"0a", X"f8", X"a6", X"05", 
    X"08", X"a6", X"06", X"08", X"a6", X"07", X"c0", X"02", 
    X"c0", X"03", X"c0", X"04", X"e5", X"0c", X"24", X"0a", 
    X"f8", X"74", X"02", X"26", X"fd", X"e4", X"08", X"36", 
    X"fe", X"08", X"86", X"07", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"70", X"5a", X"fa", X"a3", X"12", 
    X"70", X"5a", X"fb", X"a3", X"12", X"70", X"5a", X"fc", 
    X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"12", X"70", 
    X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"fb", X"e5", 
    X"0c", X"24", X"0d", X"f8", X"c3", X"e6", X"9a", X"08", 
    X"e6", X"9b", X"d0", X"04", X"d0", X"03", X"d0", X"02", 
    X"40", X"1d", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"e5", X"0c", X"24", X"0a", X"f8", X"12", X"70", X"5a", 
    X"f6", X"a3", X"12", X"70", X"5a", X"08", X"f6", X"a3", 
    X"12", X"70", X"5a", X"08", X"f6", X"80", X"97", X"e5", 
    X"0c", X"24", X"04", X"f8", X"74", X"02", X"2a", X"f6", 
    X"e4", X"3b", X"08", X"f6", X"08", X"a6", X"04", X"e5", 
    X"0c", X"24", X"0a", X"f8", X"e5", X"0c", X"24", X"07", 
    X"f9", X"74", X"02", X"26", X"f7", X"e4", X"08", X"36", 
    X"09", X"f7", X"08", X"09", X"e6", X"f7", X"e5", X"0c", 
    X"24", X"07", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"70", X"5a", X"fd", X"a3", 
    X"12", X"70", X"5a", X"fe", X"a3", X"12", X"70", X"5a", 
    X"ff", X"e5", X"0c", X"24", X"04", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"ed", X"12", 
    X"66", X"a0", X"a3", X"ee", X"12", X"66", X"a0", X"a3", 
    X"ef", X"12", X"66", X"a0", X"74", X"05", X"2d", X"fd", 
    X"e4", X"3e", X"fe", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"ea", X"12", X"66", X"a0", X"a3", X"eb", X"12", 
    X"66", X"a0", X"a3", X"ec", X"12", X"66", X"a0", X"74", 
    X"05", X"2a", X"fd", X"e4", X"3b", X"fe", X"8c", X"07", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"e5", X"0c", 
    X"24", X"0a", X"f8", X"e6", X"12", X"66", X"a0", X"a3", 
    X"08", X"e6", X"12", X"66", X"a0", X"a3", X"08", X"e6", 
    X"12", X"66", X"a0", X"e5", X"0c", X"24", X"07", X"f8", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"ea", X"12", X"66", X"a0", X"a3", X"eb", X"12", X"66", 
    X"a0", X"a3", X"ec", X"12", X"66", X"a0", X"74", X"0b", 
    X"2a", X"fa", X"e4", X"3b", X"fb", X"8a", X"82", X"8b", 
    X"83", X"8c", X"f0", X"a8", X"0c", X"08", X"e6", X"12", 
    X"66", X"a0", X"a3", X"08", X"e6", X"12", X"66", X"a0", 
    X"a3", X"08", X"e6", X"12", X"66", X"a0", X"a8", X"0c", 
    X"08", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"70", X"5a", X"ff", X"0f", X"a8", X"0c", 
    X"08", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"ef", X"12", X"66", X"a0", X"85", X"0c", X"81", 
    X"d0", X"0c", X"22", X"c0", X"0c", X"85", X"81", X"0c", 
    X"c0", X"82", X"c0", X"83", X"c0", X"f0", X"e5", X"81", 
    X"24", X"0c", X"f5", X"81", X"a8", X"0c", X"08", X"74", 
    X"0b", X"26", X"fa", X"e4", X"08", X"36", X"fb", X"08", 
    X"86", X"04", X"8a", X"82", X"8b", X"83", X"8c", X"f0", 
    X"e5", X"0c", X"24", X"0d", X"f8", X"12", X"70", X"5a", 
    X"f6", X"a3", X"12", X"70", X"5a", X"08", X"f6", X"a3", 
    X"12", X"70", X"5a", X"08", X"f6", X"a8", X"0c", X"08", 
    X"e5", X"0c", X"24", X"04", X"f9", X"74", X"02", X"26", 
    X"f7", X"e4", X"08", X"36", X"09", X"f7", X"08", X"09", 
    X"e6", X"f7", X"e5", X"0c", X"24", X"04", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"12", 
    X"70", X"5a", X"fd", X"a3", X"12", X"70", X"5a", X"fe", 
    X"a3", X"12", X"70", X"5a", X"ff", X"e5", X"0c", X"24", 
    X"0a", X"f8", X"74", X"05", X"2d", X"f6", X"e4", X"3e", 
    X"08", X"f6", X"08", X"a6", X"07", X"a8", X"0c", X"08", 
    X"e5", X"0c", X"24", X"07", X"f9", X"74", X"05", X"26", 
    X"f7", X"e4", X"08", X"36", X"09", X"f7", X"08", X"09", 
    X"e6", X"f7", X"e5", X"0c", X"24", X"07", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"12", 
    X"70", X"5a", X"fd", X"a3", X"12", X"70", X"5a", X"fe", 
    X"a3", X"12", X"70", X"5a", X"ff", X"e5", X"0c", X"24", 
    X"0a", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"ed", X"12", X"66", X"a0", X"a3", X"ee", 
    X"12", X"66", X"a0", X"a3", X"ef", X"12", X"66", X"a0", 
    X"e5", X"0c", X"24", X"07", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"fd", X"a3", X"12", X"70", X"5a", X"fe", X"a3", X"12", 
    X"70", X"5a", X"ff", X"e5", X"0c", X"24", X"0a", X"f8", 
    X"74", X"02", X"2d", X"f6", X"e4", X"3e", X"08", X"f6", 
    X"08", X"a6", X"07", X"e5", X"0c", X"24", X"04", X"f8", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"12", X"70", X"5a", X"fd", X"a3", X"12", X"70", X"5a", 
    X"fe", X"a3", X"12", X"70", X"5a", X"ff", X"e5", X"0c", 
    X"24", X"0a", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"ed", X"12", X"66", X"a0", X"a3", 
    X"ee", X"12", X"66", X"a0", X"a3", X"ef", X"12", X"66", 
    X"a0", X"e5", X"0c", X"24", X"0d", X"f8", X"e5", X"0c", 
    X"24", X"0a", X"f9", X"74", X"01", X"26", X"f7", X"e4", 
    X"08", X"36", X"09", X"f7", X"08", X"09", X"e6", X"f7", 
    X"e5", X"0c", X"24", X"0a", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"fd", X"a3", X"12", X"70", X"5a", X"fe", X"a3", X"12", 
    X"70", X"5a", X"ff", X"a8", X"0c", X"08", X"c0", X"05", 
    X"c0", X"06", X"c0", X"07", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"00", X"11", X"15", 
    X"81", X"15", X"81", X"15", X"81", X"60", X"02", X"80", 
    X"36", X"e5", X"0c", X"24", X"07", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"70", 
    X"5a", X"fd", X"a3", X"12", X"70", X"5a", X"fe", X"a3", 
    X"12", X"70", X"5a", X"ff", X"e5", X"0c", X"24", X"0a", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"ed", X"12", X"66", X"a0", X"a3", X"ee", X"12", 
    X"66", X"a0", X"a3", X"ef", X"12", X"66", X"a0", X"8a", 
    X"82", X"8b", X"83", X"8c", X"f0", X"e4", X"12", X"66", 
    X"a0", X"a3", X"12", X"66", X"a0", X"a3", X"12", X"66", 
    X"a0", X"e5", X"0c", X"24", X"0d", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"70", 
    X"5a", X"ff", X"1f", X"e5", X"0c", X"24", X"0d", X"f8", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"ef", X"12", X"66", X"a0", X"e5", X"0c", X"24", X"0d", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"70", X"5a", X"f5", X"82", X"85", X"0c", 
    X"81", X"d0", X"0c", X"22", X"c0", X"0c", X"85", X"81", 
    X"0c", X"c0", X"82", X"c0", X"83", X"c0", X"f0", X"e5", 
    X"81", X"24", X"09", X"f5", X"81", X"c0", X"e0", X"c0", 
    X"a8", X"c2", X"af", X"a8", X"0c", X"08", X"74", X"06", 
    X"26", X"fa", X"e4", X"08", X"36", X"fb", X"08", X"86", 
    X"04", X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"e5", X"0c", X"24", X"04", 
    X"f9", X"12", X"70", X"5a", X"f7", X"a3", X"12", X"70", 
    X"5a", X"09", X"f7", X"a3", X"12", X"70", X"5a", X"09", 
    X"f7", X"a8", X"0c", X"08", X"e5", X"0c", X"24", X"07", 
    X"f9", X"74", X"25", X"26", X"f7", X"e4", X"08", X"36", 
    X"09", X"f7", X"08", X"09", X"e6", X"f7", X"e5", X"0c", 
    X"24", X"07", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"70", X"5a", X"fe", X"a8", 
    X"0c", X"08", X"e5", X"0c", X"24", X"0a", X"f9", X"74", 
    X"26", X"26", X"f7", X"e4", X"08", X"36", X"09", X"f7", 
    X"08", X"09", X"e6", X"f7", X"e5", X"0c", X"24", X"0a", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"70", X"5a", X"8e", X"f0", X"a4", X"c8", 
    X"e5", X"0c", X"24", X"04", X"c8", X"26", X"fd", X"08", 
    X"e6", X"35", X"f0", X"fe", X"08", X"86", X"07", X"8a", 
    X"82", X"8b", X"83", X"8c", X"f0", X"ed", X"12", X"66", 
    X"a0", X"a3", X"ee", X"12", X"66", X"a0", X"a3", X"ef", 
    X"12", X"66", X"a0", X"a8", X"0c", X"08", X"74", X"24", 
    X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", X"86", 
    X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"e4", 
    X"12", X"66", X"a0", X"a8", X"0c", X"08", X"e5", X"0c", 
    X"24", X"04", X"f9", X"74", X"03", X"26", X"f7", X"e4", 
    X"08", X"36", X"09", X"f7", X"08", X"09", X"e6", X"f7", 
    X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"70", X"5a", X"fd", X"a3", 
    X"12", X"70", X"5a", X"fe", X"a3", X"12", X"70", X"5a", 
    X"ff", X"e5", X"0c", X"24", X"04", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"ed", X"12", 
    X"66", X"a0", X"a3", X"ee", X"12", X"66", X"a0", X"a3", 
    X"ef", X"12", X"66", X"a0", X"74", X"03", X"2a", X"fa", 
    X"e4", X"3b", X"fb", X"a8", X"0c", X"08", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"e5", X"0c", 
    X"24", X"04", X"f9", X"12", X"70", X"5a", X"f7", X"a3", 
    X"12", X"70", X"5a", X"09", X"f7", X"a3", X"12", X"70", 
    X"5a", X"09", X"f7", X"e5", X"0c", X"24", X"07", X"f8", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"12", X"70", X"5a", X"ff", X"7e", X"00", X"e5", X"0c", 
    X"24", X"07", X"f8", X"ef", X"24", X"ff", X"f6", X"ee", 
    X"34", X"ff", X"08", X"f6", X"e5", X"0c", X"24", X"0a", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"70", X"5a", X"fd", X"7f", X"00", X"c0", 
    X"04", X"c0", X"03", X"c0", X"02", X"c0", X"05", X"c0", 
    X"07", X"e5", X"0c", X"24", X"07", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"12", X"66", X"bb", X"ae", X"82", 
    X"af", X"83", X"15", X"81", X"15", X"81", X"d0", X"02", 
    X"d0", X"03", X"d0", X"04", X"e5", X"0c", X"24", X"04", 
    X"f8", X"ee", X"26", X"fe", X"ef", X"08", X"36", X"ff", 
    X"08", X"86", X"05", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"ee", X"12", X"66", X"a0", X"a3", X"ef", X"12", 
    X"66", X"a0", X"a3", X"ed", X"12", X"66", X"a0", X"a8", 
    X"0c", X"08", X"74", X"27", X"26", X"fd", X"e4", X"08", 
    X"36", X"fe", X"08", X"86", X"07", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"74", X"ff", X"12", X"66", X"a0", 
    X"a8", X"0c", X"08", X"74", X"28", X"26", X"fd", X"e4", 
    X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"74", X"ff", X"12", X"66", 
    X"a0", X"e5", X"0c", X"24", X"fd", X"f8", X"e6", X"70", 
    X"39", X"a8", X"0c", X"08", X"74", X"0c", X"26", X"fd", 
    X"e4", X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"60", X"4e", X"a8", X"0c", X"08", X"74", X"0c", X"26", 
    X"fd", X"e4", X"08", X"36", X"fe", X"08", X"86", X"07", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"10", 
    X"57", X"e5", X"82", X"60", X"33", X"12", X"64", X"b5", 
    X"80", X"2e", X"a8", X"0c", X"08", X"74", X"0c", X"26", 
    X"fd", X"e4", X"08", X"36", X"fe", X"08", X"86", X"07", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"2b", 
    X"dd", X"a8", X"0c", X"08", X"74", X"18", X"26", X"fd", 
    X"e4", X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"2b", X"dd", 
    X"d0", X"e0", X"53", X"e0", X"80", X"e5", X"e0", X"42", 
    X"a8", X"d0", X"e0", X"75", X"82", X"01", X"85", X"0c", 
    X"81", X"d0", X"0c", X"22", X"c0", X"0c", X"85", X"81", 
    X"0c", X"c0", X"82", X"e5", X"0c", X"24", X"fd", X"f8", 
    X"e6", X"70", X"04", X"fd", X"fe", X"80", X"13", X"a8", 
    X"0c", X"08", X"e5", X"0c", X"24", X"fd", X"f9", X"86", 
    X"f0", X"e7", X"a4", X"fb", X"ac", X"f0", X"8b", X"05", 
    X"8c", X"06", X"74", X"29", X"2d", X"fd", X"e4", X"3e", 
    X"fe", X"8d", X"82", X"8e", X"83", X"12", X"61", X"84", 
    X"ac", X"82", X"ad", X"83", X"ae", X"f0", X"ec", X"4d", 
    X"60", X"43", X"8c", X"02", X"8d", X"03", X"8e", X"07", 
    X"74", X"29", X"2a", X"fa", X"e4", X"3b", X"fb", X"c0", 
    X"06", X"c0", X"05", X"c0", X"04", X"c0", X"04", X"c0", 
    X"05", X"c0", X"06", X"e5", X"0c", X"24", X"fc", X"f8", 
    X"e6", X"c0", X"e0", X"c0", X"02", X"c0", X"03", X"c0", 
    X"07", X"e5", X"0c", X"24", X"fd", X"f8", X"e6", X"c0", 
    X"e0", X"a8", X"0c", X"08", X"86", X"82", X"12", X"35", 
    X"30", X"e5", X"81", X"24", X"f8", X"f5", X"81", X"d0", 
    X"04", X"d0", X"05", X"d0", X"06", X"8c", X"82", X"8d", 
    X"83", X"8e", X"f0", X"15", X"81", X"d0", X"0c", X"22", 
    X"c0", X"0c", X"85", X"81", X"0c", X"c0", X"82", X"e5", 
    X"0c", X"24", X"fd", X"f8", X"e6", X"70", X"30", X"e5", 
    X"0c", X"24", X"f6", X"f8", X"86", X"04", X"08", X"86", 
    X"05", X"08", X"86", X"06", X"e5", X"0c", X"24", X"f6", 
    X"f8", X"86", X"02", X"08", X"86", X"03", X"08", X"86", 
    X"07", X"8c", X"82", X"8d", X"83", X"8e", X"f0", X"ea", 
    X"12", X"66", X"a0", X"a3", X"eb", X"12", X"66", X"a0", 
    X"a3", X"ef", X"12", X"66", X"a0", X"80", X"2e", X"e5", 
    X"0c", X"24", X"f6", X"f8", X"86", X"04", X"08", X"86", 
    X"05", X"08", X"86", X"06", X"e5", X"0c", X"24", X"fa", 
    X"f8", X"86", X"02", X"08", X"86", X"03", X"08", X"86", 
    X"07", X"8c", X"82", X"8d", X"83", X"8e", X"f0", X"ea", 
    X"12", X"66", X"a0", X"a3", X"eb", X"12", X"66", X"a0", 
    X"a3", X"ef", X"12", X"66", X"a0", X"e5", X"0c", X"24", 
    X"f6", X"f8", X"86", X"05", X"08", X"86", X"06", X"08", 
    X"86", X"07", X"74", X"25", X"2d", X"fa", X"e4", X"3e", 
    X"fb", X"8f", X"04", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"a8", X"0c", X"08", X"e6", X"12", X"66", X"a0", 
    X"74", X"26", X"2d", X"fa", X"e4", X"3e", X"fb", X"8f", 
    X"04", X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"e5", 
    X"0c", X"24", X"fd", X"f8", X"e6", X"12", X"66", X"a0", 
    X"74", X"01", X"c0", X"e0", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"32", X"34", X"15", X"81", X"15", 
    X"81", X"d0", X"0c", X"22", X"c0", X"0c", X"e5", X"81", 
    X"f5", X"0c", X"24", X"11", X"f5", X"81", X"ad", X"82", 
    X"ab", X"83", X"ac", X"f0", X"e5", X"0c", X"24", X"0b", 
    X"f8", X"76", X"00", X"e5", X"0c", X"24", X"0f", X"f8", 
    X"a6", X"05", X"08", X"a6", X"03", X"08", X"a6", X"04", 
    X"e5", X"0c", X"24", X"f8", X"f8", X"e4", X"b6", X"02", 
    X"01", X"04", X"ff", X"e5", X"0c", X"24", X"0c", X"fe", 
    X"e5", X"0c", X"24", X"07", X"f8", X"a6", X"06", X"a8", 
    X"0c", X"08", X"74", X"24", X"2d", X"f6", X"e4", X"3b", 
    X"08", X"f6", X"08", X"a6", X"04", X"e5", X"0c", X"24", 
    X"04", X"f8", X"74", X"25", X"2d", X"f6", X"e4", X"3b", 
    X"08", X"f6", X"08", X"a6", X"04", X"c0", X"e0", X"c0", 
    X"a8", X"c2", X"af", X"a8", X"0c", X"08", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"70", 
    X"5a", X"fd", X"e5", X"0c", X"24", X"04", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"12", 
    X"70", X"5a", X"fc", X"c3", X"ed", X"9c", X"40", X"06", 
    X"ef", X"70", X"03", X"02", X"36", X"fc", X"e5", X"0c", 
    X"24", X"f8", X"f8", X"e6", X"c0", X"e0", X"e5", X"0c", 
    X"24", X"fb", X"f8", X"e6", X"c0", X"e0", X"08", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"e5", X"0c", 
    X"24", X"0f", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"44", X"bd", X"ac", X"82", 
    X"e5", X"81", X"24", X"fc", X"f5", X"81", X"8c", X"07", 
    X"e5", X"0c", X"24", X"0f", X"f8", X"74", X"18", X"26", 
    X"fa", X"e4", X"08", X"36", X"fb", X"08", X"86", X"04", 
    X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"12", X"70", 
    X"5a", X"60", X"22", X"e5", X"0c", X"24", X"0f", X"f8", 
    X"74", X"18", X"26", X"fa", X"e4", X"08", X"36", X"fb", 
    X"08", X"86", X"04", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"12", X"10", X"57", X"e5", X"82", X"60", X"0b", 
    X"12", X"64", X"b5", X"80", X"06", X"ef", X"60", X"03", 
    X"12", X"64", X"b5", X"d0", X"e0", X"53", X"e0", X"80", 
    X"e5", X"e0", X"42", X"a8", X"d0", X"e0", X"75", X"82", 
    X"01", X"02", X"38", X"9e", X"e5", X"0c", X"24", X"f9", 
    X"f8", X"e6", X"08", X"46", X"70", X"11", X"d0", X"e0", 
    X"53", X"e0", X"80", X"e5", X"e0", X"42", X"a8", X"d0", 
    X"e0", X"75", X"82", X"00", X"02", X"38", X"9e", X"e5", 
    X"0c", X"24", X"0b", X"f8", X"e6", X"70", X"1d", X"8e", 
    X"02", X"fb", X"7c", X"40", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"c0", X"07", X"c0", X"06", X"12", X"13", 
    X"1e", X"d0", X"06", X"d0", X"07", X"e5", X"0c", X"24", 
    X"0b", X"f8", X"76", X"01", X"d0", X"e0", X"53", X"e0", 
    X"80", X"e5", X"e0", X"42", X"a8", X"d0", X"e0", X"c0", 
    X"07", X"c0", X"06", X"12", X"09", X"4a", X"d0", X"06", 
    X"d0", X"07", X"c0", X"e0", X"c0", X"a8", X"c2", X"af", 
    X"e5", X"0c", X"24", X"0f", X"f8", X"74", X"27", X"26", 
    X"fa", X"e4", X"08", X"36", X"fb", X"08", X"86", X"04", 
    X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"12", X"70", 
    X"5a", X"fd", X"bd", X"ff", X"0a", X"8a", X"82", X"8b", 
    X"83", X"8c", X"f0", X"e4", X"12", X"66", X"a0", X"e5", 
    X"0c", X"24", X"0f", X"f8", X"74", X"28", X"26", X"fa", 
    X"e4", X"08", X"36", X"fb", X"08", X"86", X"04", X"8a", 
    X"82", X"8b", X"83", X"8c", X"f0", X"12", X"70", X"5a", 
    X"fd", X"bd", X"ff", X"0a", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"e4", X"12", X"66", X"a0", X"c0", X"07", 
    X"d0", X"e0", X"53", X"e0", X"80", X"e5", X"e0", X"42", 
    X"a8", X"d0", X"e0", X"e5", X"0c", X"24", X"f9", X"fc", 
    X"e5", X"0c", X"24", X"08", X"f8", X"a6", X"04", X"08", 
    X"76", X"00", X"08", X"76", X"40", X"e5", X"0c", X"24", 
    X"07", X"f8", X"86", X"04", X"7d", X"00", X"7f", X"40", 
    X"c0", X"06", X"e5", X"0c", X"24", X"08", X"f8", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"08", X"e6", 
    X"c0", X"e0", X"8c", X"82", X"8d", X"83", X"8f", X"f0", 
    X"12", X"13", X"4e", X"af", X"82", X"15", X"81", X"15", 
    X"81", X"15", X"81", X"d0", X"06", X"ef", X"d0", X"07", 
    X"60", X"03", X"02", X"38", X"88", X"e5", X"0c", X"24", 
    X"0f", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"c0", X"07", X"c0", X"06", X"12", X"4b", 
    X"1f", X"e5", X"82", X"d0", X"06", X"d0", X"07", X"60", 
    X"51", X"e5", X"0c", X"24", X"0f", X"f8", X"74", X"0c", 
    X"26", X"fb", X"e4", X"08", X"36", X"fc", X"08", X"86", 
    X"05", X"c0", X"07", X"c0", X"06", X"e5", X"0c", X"24", 
    X"f9", X"f8", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"8b", X"82", X"8c", X"83", X"8d", X"f0", X"12", 
    X"0f", X"92", X"15", X"81", X"15", X"81", X"e5", X"0c", 
    X"24", X"0f", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"49", X"52", X"12", X"09", 
    X"52", X"e5", X"82", X"d0", X"06", X"d0", X"07", X"60", 
    X"03", X"02", X"36", X"45", X"12", X"64", X"b5", X"02", 
    X"36", X"45", X"e5", X"0c", X"24", X"0f", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"c0", 
    X"07", X"c0", X"06", X"12", X"49", X"52", X"12", X"09", 
    X"52", X"d0", X"06", X"d0", X"07", X"02", X"36", X"45", 
    X"e5", X"0c", X"24", X"0f", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"49", X"52", 
    X"12", X"09", X"52", X"75", X"82", X"00", X"85", X"0c", 
    X"81", X"d0", X"0c", X"22", X"c0", X"0c", X"85", X"81", 
    X"0c", X"05", X"81", X"05", X"81", X"05", X"81", X"aa", 
    X"82", X"ab", X"83", X"ac", X"f0", X"a8", X"0c", X"08", 
    X"a6", X"02", X"08", X"a6", X"03", X"08", X"a6", X"04", 
    X"74", X"24", X"2a", X"fd", X"e4", X"3b", X"fe", X"8c", 
    X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"70", X"5a", X"fd", X"74", X"25", X"2a", X"fc", X"e4", 
    X"3b", X"fe", X"8c", X"07", X"8c", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"70", X"5a", X"fc", X"c3", X"ed", 
    X"9c", X"40", X"0d", X"e5", X"0c", X"24", X"f7", X"f8", 
    X"b6", X"02", X"02", X"80", X"03", X"02", X"39", X"b9", 
    X"a8", X"0c", X"08", X"74", X"28", X"26", X"fd", X"e4", 
    X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"ff", 
    X"c0", X"07", X"e5", X"0c", X"24", X"f7", X"f8", X"e6", 
    X"c0", X"e0", X"e5", X"0c", X"24", X"fb", X"f8", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"08", X"e6", 
    X"c0", X"e0", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"44", X"bd", 
    X"e5", X"81", X"24", X"fc", X"f5", X"81", X"d0", X"07", 
    X"bf", X"ff", X"58", X"a8", X"0c", X"08", X"74", X"18", 
    X"26", X"fc", X"e4", X"08", X"36", X"fd", X"08", X"86", 
    X"06", X"8c", X"82", X"8d", X"83", X"8e", X"f0", X"12", 
    X"70", X"5a", X"60", X"58", X"a8", X"0c", X"08", X"74", 
    X"18", X"26", X"fc", X"e4", X"08", X"36", X"fd", X"08", 
    X"86", X"06", X"8c", X"82", X"8d", X"83", X"8e", X"f0", 
    X"12", X"10", X"57", X"e5", X"82", X"60", X"3d", X"e5", 
    X"0c", X"24", X"f8", X"f8", X"e6", X"08", X"46", X"60", 
    X"33", X"e5", X"0c", X"24", X"f8", X"f8", X"86", X"04", 
    X"08", X"86", X"05", X"08", X"86", X"06", X"8c", X"82", 
    X"8d", X"83", X"8e", X"f0", X"74", X"01", X"12", X"66", 
    X"a0", X"80", X"19", X"a8", X"0c", X"08", X"74", X"28", 
    X"26", X"fc", X"e4", X"08", X"36", X"fd", X"08", X"86", 
    X"06", X"0f", X"8c", X"82", X"8d", X"83", X"8e", X"f0", 
    X"ef", X"12", X"66", X"a0", X"75", X"82", X"01", X"80", 
    X"03", X"75", X"82", X"00", X"85", X"0c", X"81", X"d0", 
    X"0c", X"22", X"c0", X"0c", X"85", X"81", X"0c", X"c0", 
    X"82", X"c0", X"83", X"c0", X"f0", X"e5", X"81", X"24", 
    X"04", X"f5", X"81", X"a8", X"0c", X"08", X"74", X"24", 
    X"26", X"fa", X"e4", X"08", X"36", X"fb", X"08", X"86", 
    X"04", X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"e5", 
    X"0c", X"24", X"07", X"f8", X"12", X"70", X"5a", X"f6", 
    X"a8", X"0c", X"08", X"74", X"25", X"26", X"fd", X"e4", 
    X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fd", 
    X"e5", X"0c", X"24", X"07", X"f8", X"c3", X"e6", X"9d", 
    X"40", X"03", X"02", X"3a", X"be", X"a8", X"0c", X"08", 
    X"e5", X"0c", X"24", X"04", X"f9", X"74", X"28", X"26", 
    X"f7", X"e4", X"08", X"36", X"09", X"f7", X"08", X"09", 
    X"e6", X"f7", X"e5", X"0c", X"24", X"04", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"12", 
    X"70", X"5a", X"ff", X"e5", X"0c", X"24", X"07", X"f8", 
    X"e6", X"04", X"fe", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"12", X"66", X"a0", X"bf", X"ff", X"58", X"a8", 
    X"0c", X"08", X"74", X"18", X"26", X"fc", X"e4", X"08", 
    X"36", X"fd", X"08", X"86", X"06", X"8c", X"82", X"8d", 
    X"83", X"8e", X"f0", X"12", X"70", X"5a", X"60", X"51", 
    X"a8", X"0c", X"08", X"74", X"18", X"26", X"fc", X"e4", 
    X"08", X"36", X"fd", X"08", X"86", X"06", X"8c", X"82", 
    X"8d", X"83", X"8e", X"f0", X"12", X"10", X"57", X"e5", 
    X"82", X"60", X"36", X"e5", X"0c", X"24", X"fb", X"f8", 
    X"e6", X"08", X"46", X"60", X"2c", X"e5", X"0c", X"24", 
    X"fb", X"f8", X"86", X"04", X"08", X"86", X"05", X"08", 
    X"86", X"06", X"8c", X"82", X"8d", X"83", X"8e", X"f0", 
    X"74", X"01", X"12", X"66", X"a0", X"80", X"12", X"0f", 
    X"e5", X"0c", X"24", X"04", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"ef", X"12", X"66", 
    X"a0", X"75", X"82", X"01", X"80", X"03", X"75", X"82", 
    X"00", X"85", X"0c", X"81", X"d0", X"0c", X"22", X"c0", 
    X"0c", X"e5", X"81", X"f5", X"0c", X"24", X"0b", X"f5", 
    X"81", X"ac", X"82", X"ad", X"83", X"af", X"f0", X"e5", 
    X"0c", X"24", X"05", X"f8", X"76", X"00", X"e5", X"0c", 
    X"24", X"09", X"f8", X"a6", X"04", X"08", X"a6", X"05", 
    X"08", X"a6", X"07", X"e5", X"0c", X"24", X"06", X"fe", 
    X"e5", X"0c", X"24", X"04", X"f8", X"a6", X"06", X"a8", 
    X"0c", X"08", X"74", X"24", X"2c", X"f6", X"e4", X"3d", 
    X"08", X"f6", X"08", X"a6", X"07", X"c0", X"e0", X"c0", 
    X"a8", X"c2", X"af", X"a8", X"0c", X"08", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"70", 
    X"5a", X"fc", X"fd", X"70", X"03", X"02", X"3b", X"b2", 
    X"c0", X"05", X"e5", X"0c", X"24", X"fb", X"f8", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"08", X"e6", 
    X"c0", X"e0", X"e5", X"0c", X"24", X"09", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"12", 
    X"48", X"02", X"15", X"81", X"15", X"81", X"15", X"81", 
    X"d0", X"05", X"e5", X"0c", X"24", X"09", X"f8", X"74", 
    X"24", X"26", X"fb", X"e4", X"08", X"36", X"fc", X"08", 
    X"86", X"07", X"ed", X"14", X"fa", X"8b", X"82", X"8c", 
    X"83", X"8f", X"f0", X"12", X"66", X"a0", X"e5", X"0c", 
    X"24", X"09", X"f8", X"74", X"0c", X"26", X"fb", X"e4", 
    X"08", X"36", X"fc", X"08", X"86", X"07", X"8b", X"82", 
    X"8c", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"60", 
    X"20", X"e5", X"0c", X"24", X"09", X"f8", X"74", X"0c", 
    X"26", X"fb", X"e4", X"08", X"36", X"fc", X"08", X"86", 
    X"07", X"8b", X"82", X"8c", X"83", X"8f", X"f0", X"12", 
    X"10", X"57", X"e5", X"82", X"60", X"03", X"12", X"64", 
    X"b5", X"d0", X"e0", X"53", X"e0", X"80", X"e5", X"e0", 
    X"42", X"a8", X"d0", X"e0", X"75", X"82", X"01", X"02", 
    X"3d", X"48", X"e5", X"0c", X"24", X"f9", X"f8", X"e6", 
    X"08", X"46", X"70", X"11", X"d0", X"e0", X"53", X"e0", 
    X"80", X"e5", X"e0", X"42", X"a8", X"d0", X"e0", X"75", 
    X"82", X"00", X"02", X"3d", X"48", X"e5", X"0c", X"24", 
    X"05", X"f8", X"e6", X"70", X"19", X"8e", X"03", X"fc", 
    X"7f", X"40", X"8b", X"82", X"8c", X"83", X"8f", X"f0", 
    X"c0", X"06", X"12", X"13", X"1e", X"d0", X"06", X"e5", 
    X"0c", X"24", X"05", X"f8", X"76", X"01", X"d0", X"e0", 
    X"53", X"e0", X"80", X"e5", X"e0", X"42", X"a8", X"d0", 
    X"e0", X"c0", X"06", X"12", X"09", X"4a", X"d0", X"06", 
    X"c0", X"e0", X"c0", X"a8", X"c2", X"af", X"e5", X"0c", 
    X"24", X"09", X"f8", X"74", X"27", X"26", X"fb", X"e4", 
    X"08", X"36", X"fc", X"08", X"86", X"07", X"8b", X"82", 
    X"8c", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fa", 
    X"ba", X"ff", X"0a", X"8b", X"82", X"8c", X"83", X"8f", 
    X"f0", X"e4", X"12", X"66", X"a0", X"e5", X"0c", X"24", 
    X"09", X"f8", X"74", X"28", X"26", X"fb", X"e4", X"08", 
    X"36", X"fc", X"08", X"86", X"07", X"8b", X"82", X"8c", 
    X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fa", X"ba", 
    X"ff", X"0a", X"8b", X"82", X"8c", X"83", X"8f", X"f0", 
    X"e4", X"12", X"66", X"a0", X"c0", X"06", X"d0", X"e0", 
    X"53", X"e0", X"80", X"e5", X"e0", X"42", X"a8", X"d0", 
    X"e0", X"e5", X"0c", X"24", X"f9", X"ff", X"7c", X"00", 
    X"7b", X"40", X"e5", X"0c", X"24", X"04", X"f8", X"86", 
    X"02", X"7d", X"00", X"7e", X"40", X"c0", X"06", X"c0", 
    X"07", X"c0", X"04", X"c0", X"03", X"8a", X"82", X"8d", 
    X"83", X"8e", X"f0", X"12", X"13", X"4e", X"af", X"82", 
    X"15", X"81", X"15", X"81", X"15", X"81", X"d0", X"06", 
    X"d0", X"06", X"ef", X"60", X"03", X"02", X"3d", X"17", 
    X"e5", X"0c", X"24", X"09", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"c0", X"06", X"12", 
    X"4a", X"cc", X"e5", X"82", X"d0", X"06", X"60", X"4d", 
    X"e5", X"0c", X"24", X"09", X"f8", X"74", X"18", X"26", 
    X"fc", X"e4", X"08", X"36", X"fd", X"08", X"86", X"07", 
    X"c0", X"06", X"e5", X"0c", X"24", X"f9", X"f8", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"8c", X"82", 
    X"8d", X"83", X"8f", X"f0", X"12", X"0f", X"92", X"15", 
    X"81", X"15", X"81", X"e5", X"0c", X"24", X"09", X"f8", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"12", X"49", X"52", X"12", X"09", X"52", X"e5", X"82", 
    X"d0", X"06", X"60", X"03", X"02", X"3b", X"05", X"12", 
    X"64", X"b5", X"02", X"3b", X"05", X"e5", X"0c", X"24", 
    X"09", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"c0", X"06", X"12", X"49", X"52", X"12", 
    X"09", X"52", X"d0", X"06", X"02", X"3b", X"05", X"e5", 
    X"0c", X"24", X"09", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"c0", X"06", X"12", X"49", 
    X"52", X"12", X"09", X"52", X"e5", X"0c", X"24", X"09", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"4a", X"cc", X"e5", X"82", X"d0", X"06", 
    X"70", X"03", X"02", X"3b", X"05", X"75", X"82", X"00", 
    X"85", X"0c", X"81", X"d0", X"0c", X"22", X"c0", X"0c", 
    X"e5", X"81", X"f5", X"0c", X"24", X"0b", X"f5", X"81", 
    X"ac", X"82", X"ad", X"83", X"af", X"f0", X"e5", X"0c", 
    X"24", X"0b", X"f8", X"76", X"00", X"e5", X"0c", X"24", 
    X"08", X"f8", X"a6", X"04", X"08", X"a6", X"05", X"08", 
    X"a6", X"07", X"e5", X"0c", X"24", X"05", X"fe", X"e5", 
    X"0c", X"24", X"04", X"f8", X"a6", X"06", X"a8", X"0c", 
    X"08", X"74", X"24", X"2c", X"f6", X"e4", X"3d", X"08", 
    X"f6", X"08", X"a6", X"07", X"c0", X"e0", X"c0", X"a8", 
    X"c2", X"af", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"fc", X"ff", X"60", X"5e", X"ef", X"14", X"fc", X"a8", 
    X"0c", X"08", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"ec", X"12", X"66", X"a0", X"e5", X"0c", 
    X"24", X"08", X"f8", X"74", X"0c", X"26", X"fb", X"e4", 
    X"08", X"36", X"fc", X"08", X"86", X"07", X"8b", X"82", 
    X"8c", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"60", 
    X"20", X"e5", X"0c", X"24", X"08", X"f8", X"74", X"0c", 
    X"26", X"fb", X"e4", X"08", X"36", X"fc", X"08", X"86", 
    X"07", X"8b", X"82", X"8c", X"83", X"8f", X"f0", X"12", 
    X"10", X"57", X"e5", X"82", X"60", X"03", X"12", X"64", 
    X"b5", X"d0", X"e0", X"53", X"e0", X"80", X"e5", X"e0", 
    X"42", X"a8", X"d0", X"e0", X"75", X"82", X"01", X"02", 
    X"3f", X"98", X"e5", X"0c", X"24", X"fc", X"f8", X"e6", 
    X"08", X"46", X"70", X"11", X"d0", X"e0", X"53", X"e0", 
    X"80", X"e5", X"e0", X"42", X"a8", X"d0", X"e0", X"75", 
    X"82", X"00", X"02", X"3f", X"98", X"e5", X"0c", X"24", 
    X"0b", X"f8", X"e6", X"70", X"19", X"8e", X"03", X"fc", 
    X"7f", X"40", X"8b", X"82", X"8c", X"83", X"8f", X"f0", 
    X"c0", X"06", X"12", X"13", X"1e", X"d0", X"06", X"e5", 
    X"0c", X"24", X"0b", X"f8", X"76", X"01", X"d0", X"e0", 
    X"53", X"e0", X"80", X"e5", X"e0", X"42", X"a8", X"d0", 
    X"e0", X"c0", X"06", X"12", X"09", X"4a", X"d0", X"06", 
    X"c0", X"e0", X"c0", X"a8", X"c2", X"af", X"e5", X"0c", 
    X"24", X"08", X"f8", X"74", X"27", X"26", X"fb", X"e4", 
    X"08", X"36", X"fc", X"08", X"86", X"07", X"8b", X"82", 
    X"8c", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fa", 
    X"ba", X"ff", X"0a", X"8b", X"82", X"8c", X"83", X"8f", 
    X"f0", X"e4", X"12", X"66", X"a0", X"e5", X"0c", X"24", 
    X"08", X"f8", X"74", X"28", X"26", X"fb", X"e4", X"08", 
    X"36", X"fc", X"08", X"86", X"07", X"8b", X"82", X"8c", 
    X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fa", X"ba", 
    X"ff", X"0a", X"8b", X"82", X"8c", X"83", X"8f", X"f0", 
    X"e4", X"12", X"66", X"a0", X"c0", X"06", X"d0", X"e0", 
    X"53", X"e0", X"80", X"e5", X"e0", X"42", X"a8", X"d0", 
    X"e0", X"e5", X"0c", X"24", X"fc", X"ff", X"7c", X"00", 
    X"7b", X"40", X"e5", X"0c", X"24", X"04", X"f8", X"86", 
    X"02", X"7d", X"00", X"7e", X"40", X"c0", X"06", X"c0", 
    X"07", X"c0", X"04", X"c0", X"03", X"8a", X"82", X"8d", 
    X"83", X"8e", X"f0", X"12", X"13", X"4e", X"af", X"82", 
    X"15", X"81", X"15", X"81", X"15", X"81", X"d0", X"06", 
    X"d0", X"06", X"ef", X"60", X"03", X"02", X"3f", X"67", 
    X"e5", X"0c", X"24", X"08", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"c0", X"06", X"12", 
    X"4a", X"cc", X"e5", X"82", X"d0", X"06", X"60", X"4d", 
    X"e5", X"0c", X"24", X"08", X"f8", X"74", X"18", X"26", 
    X"fc", X"e4", X"08", X"36", X"fd", X"08", X"86", X"07", 
    X"c0", X"06", X"e5", X"0c", X"24", X"fc", X"f8", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"8c", X"82", 
    X"8d", X"83", X"8f", X"f0", X"12", X"0f", X"92", X"15", 
    X"81", X"15", X"81", X"e5", X"0c", X"24", X"08", X"f8", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"12", X"49", X"52", X"12", X"09", X"52", X"e5", X"82", 
    X"d0", X"06", X"60", X"03", X"02", X"3d", X"8c", X"12", 
    X"64", X"b5", X"02", X"3d", X"8c", X"e5", X"0c", X"24", 
    X"08", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"c0", X"06", X"12", X"49", X"52", X"12", 
    X"09", X"52", X"d0", X"06", X"02", X"3d", X"8c", X"e5", 
    X"0c", X"24", X"08", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"c0", X"06", X"12", X"49", 
    X"52", X"12", X"09", X"52", X"e5", X"0c", X"24", X"08", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"4a", X"cc", X"e5", X"82", X"d0", X"06", 
    X"70", X"03", X"02", X"3d", X"8c", X"75", X"82", X"00", 
    X"85", X"0c", X"81", X"d0", X"0c", X"22", X"c0", X"0c", 
    X"e5", X"81", X"f5", X"0c", X"24", X"0d", X"f5", X"81", 
    X"ad", X"82", X"ab", X"83", X"af", X"f0", X"7c", X"00", 
    X"e5", X"0c", X"24", X"0b", X"f8", X"a6", X"05", X"08", 
    X"a6", X"03", X"08", X"a6", X"07", X"e5", X"0c", X"24", 
    X"08", X"fe", X"e5", X"0c", X"24", X"04", X"f8", X"a6", 
    X"06", X"a8", X"0c", X"08", X"74", X"24", X"2d", X"f6", 
    X"e4", X"3b", X"08", X"f6", X"08", X"a6", X"07", X"c0", 
    X"e0", X"c0", X"a8", X"c2", X"af", X"a8", X"0c", X"08", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"12", X"70", X"5a", X"70", X"03", X"02", X"40", X"c4", 
    X"e5", X"0c", X"24", X"0b", X"f8", X"74", X"06", X"26", 
    X"fa", X"e4", X"08", X"36", X"fb", X"08", X"86", X"07", 
    X"74", X"03", X"2a", X"fa", X"e4", X"3b", X"fb", X"8a", 
    X"82", X"8b", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"fe", X"a3", X"12", X"70", X"5a", X"fd", X"a3", X"12", 
    X"70", X"5a", X"fc", X"c0", X"06", X"c0", X"05", X"c0", 
    X"04", X"e5", X"0c", X"24", X"fb", X"f8", X"e6", X"c0", 
    X"e0", X"08", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"e5", X"0c", X"24", X"0b", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"48", 
    X"02", X"15", X"81", X"15", X"81", X"15", X"81", X"d0", 
    X"04", X"d0", X"05", X"d0", X"06", X"e5", X"0c", X"24", 
    X"0b", X"f8", X"74", X"06", X"26", X"fa", X"e4", X"08", 
    X"36", X"fb", X"08", X"86", X"07", X"74", X"03", X"2a", 
    X"fa", X"e4", X"3b", X"fb", X"8a", X"82", X"8b", X"83", 
    X"8f", X"f0", X"ee", X"12", X"66", X"a0", X"a3", X"ed", 
    X"12", X"66", X"a0", X"a3", X"ec", X"12", X"66", X"a0", 
    X"e5", X"0c", X"24", X"0b", X"f8", X"74", X"18", X"26", 
    X"fa", X"e4", X"08", X"36", X"fb", X"08", X"86", X"07", 
    X"8a", X"82", X"8b", X"83", X"8f", X"f0", X"12", X"70", 
    X"5a", X"60", X"20", X"e5", X"0c", X"24", X"0b", X"f8", 
    X"74", X"18", X"26", X"fa", X"e4", X"08", X"36", X"fb", 
    X"08", X"86", X"07", X"8a", X"82", X"8b", X"83", X"8f", 
    X"f0", X"12", X"10", X"57", X"e5", X"82", X"60", X"03", 
    X"12", X"64", X"b5", X"d0", X"e0", X"53", X"e0", X"80", 
    X"e5", X"e0", X"42", X"a8", X"d0", X"e0", X"75", X"82", 
    X"01", X"02", X"42", X"7b", X"e5", X"0c", X"24", X"f9", 
    X"f8", X"e6", X"08", X"46", X"70", X"11", X"d0", X"e0", 
    X"53", X"e0", X"80", X"e5", X"e0", X"42", X"a8", X"d0", 
    X"e0", X"75", X"82", X"00", X"02", X"42", X"7b", X"ec", 
    X"70", X"14", X"8e", X"02", X"fb", X"7f", X"40", X"8a", 
    X"82", X"8b", X"83", X"8f", X"f0", X"c0", X"06", X"12", 
    X"13", X"1e", X"d0", X"06", X"7c", X"01", X"d0", X"e0", 
    X"53", X"e0", X"80", X"e5", X"e0", X"42", X"a8", X"d0", 
    X"e0", X"c0", X"06", X"c0", X"04", X"12", X"09", X"4a", 
    X"d0", X"04", X"d0", X"06", X"c0", X"e0", X"c0", X"a8", 
    X"c2", X"af", X"e5", X"0c", X"24", X"0b", X"f8", X"74", 
    X"27", X"26", X"fa", X"e4", X"08", X"36", X"fb", X"08", 
    X"86", X"07", X"8a", X"82", X"8b", X"83", X"8f", X"f0", 
    X"12", X"70", X"5a", X"fd", X"bd", X"ff", X"0a", X"8a", 
    X"82", X"8b", X"83", X"8f", X"f0", X"e4", X"12", X"66", 
    X"a0", X"e5", X"0c", X"24", X"0b", X"f8", X"74", X"28", 
    X"26", X"fa", X"e4", X"08", X"36", X"fb", X"08", X"86", 
    X"07", X"8a", X"82", X"8b", X"83", X"8f", X"f0", X"12", 
    X"70", X"5a", X"fd", X"bd", X"ff", X"0a", X"8a", X"82", 
    X"8b", X"83", X"8f", X"f0", X"e4", X"12", X"66", X"a0", 
    X"c0", X"04", X"d0", X"e0", X"53", X"e0", X"80", X"e5", 
    X"e0", X"42", X"a8", X"d0", X"e0", X"e5", X"0c", X"24", 
    X"f9", X"ff", X"e5", X"0c", X"24", X"05", X"f8", X"a6", 
    X"07", X"08", X"76", X"00", X"08", X"76", X"40", X"e5", 
    X"0c", X"24", X"04", X"f8", X"86", X"04", X"7d", X"00", 
    X"7f", X"40", X"c0", X"06", X"c0", X"04", X"e5", X"0c", 
    X"24", X"05", X"f8", X"e6", X"c0", X"e0", X"08", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"8c", X"82", 
    X"8d", X"83", X"8f", X"f0", X"12", X"13", X"4e", X"af", 
    X"82", X"15", X"81", X"15", X"81", X"15", X"81", X"d0", 
    X"04", X"d0", X"06", X"d0", X"04", X"ef", X"60", X"03", 
    X"02", X"42", X"46", X"e5", X"0c", X"24", X"0b", X"f8", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"c0", X"06", X"c0", X"04", X"12", X"4a", X"cc", X"e5", 
    X"82", X"d0", X"04", X"d0", X"06", X"60", X"51", X"e5", 
    X"0c", X"24", X"0b", X"f8", X"74", X"18", X"26", X"fb", 
    X"e4", X"08", X"36", X"fd", X"08", X"86", X"07", X"c0", 
    X"06", X"c0", X"04", X"e5", X"0c", X"24", X"f9", X"f8", 
    X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"8b", 
    X"82", X"8d", X"83", X"8f", X"f0", X"12", X"0f", X"92", 
    X"15", X"81", X"15", X"81", X"e5", X"0c", X"24", X"0b", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"49", X"52", X"12", X"09", X"52", X"e5", 
    X"82", X"d0", X"04", X"d0", X"06", X"60", X"03", X"02", 
    X"3f", X"d7", X"12", X"64", X"b5", X"02", X"3f", X"d7", 
    X"e5", X"0c", X"24", X"0b", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"c0", X"06", X"c0", 
    X"04", X"12", X"49", X"52", X"12", X"09", X"52", X"d0", 
    X"04", X"d0", X"06", X"02", X"3f", X"d7", X"e5", X"0c", 
    X"24", X"0b", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"c0", X"06", X"c0", X"04", X"12", 
    X"49", X"52", X"12", X"09", X"52", X"e5", X"0c", X"24", 
    X"0b", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"12", X"4a", X"cc", X"e5", X"82", X"d0", 
    X"04", X"d0", X"06", X"70", X"03", X"02", X"3f", X"d7", 
    X"75", X"82", X"00", X"85", X"0c", X"81", X"d0", X"0c", 
    X"22", X"c0", X"0c", X"85", X"81", X"0c", X"c0", X"82", 
    X"c0", X"83", X"c0", X"f0", X"a8", X"0c", X"08", X"74", 
    X"24", X"26", X"fa", X"e4", X"08", X"36", X"fb", X"08", 
    X"86", X"04", X"8a", X"82", X"8b", X"83", X"8c", X"f0", 
    X"12", X"70", X"5a", X"fa", X"fc", X"70", X"03", X"02", 
    X"43", X"80", X"a8", X"0c", X"08", X"74", X"27", X"26", 
    X"fa", X"e4", X"08", X"36", X"fb", X"08", X"86", X"07", 
    X"8a", X"82", X"8b", X"83", X"8f", X"f0", X"12", X"70", 
    X"5a", X"ff", X"c0", X"07", X"c0", X"04", X"e5", X"0c", 
    X"24", X"fb", X"f8", X"e6", X"c0", X"e0", X"08", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"a8", X"0c", 
    X"08", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"48", X"02", X"15", X"81", X"15", X"81", 
    X"15", X"81", X"d0", X"04", X"d0", X"07", X"a8", X"0c", 
    X"08", X"74", X"24", X"26", X"fb", X"e4", X"08", X"36", 
    X"fd", X"08", X"86", X"06", X"1c", X"8b", X"82", X"8d", 
    X"83", X"8e", X"f0", X"ec", X"12", X"66", X"a0", X"bf", 
    X"ff", X"58", X"a8", X"0c", X"08", X"74", X"0c", X"26", 
    X"fc", X"e4", X"08", X"36", X"fd", X"08", X"86", X"06", 
    X"8c", X"82", X"8d", X"83", X"8e", X"f0", X"12", X"70", 
    X"5a", X"60", X"58", X"a8", X"0c", X"08", X"74", X"0c", 
    X"26", X"fc", X"e4", X"08", X"36", X"fd", X"08", X"86", 
    X"06", X"8c", X"82", X"8d", X"83", X"8e", X"f0", X"12", 
    X"10", X"57", X"e5", X"82", X"60", X"3d", X"e5", X"0c", 
    X"24", X"f8", X"f8", X"e6", X"08", X"46", X"60", X"33", 
    X"e5", X"0c", X"24", X"f8", X"f8", X"86", X"04", X"08", 
    X"86", X"05", X"08", X"86", X"06", X"8c", X"82", X"8d", 
    X"83", X"8e", X"f0", X"74", X"01", X"12", X"66", X"a0", 
    X"80", X"19", X"a8", X"0c", X"08", X"74", X"27", X"26", 
    X"fc", X"e4", X"08", X"36", X"fd", X"08", X"86", X"06", 
    X"0f", X"8c", X"82", X"8d", X"83", X"8e", X"f0", X"ef", 
    X"12", X"66", X"a0", X"75", X"82", X"01", X"80", X"03", 
    X"75", X"82", X"00", X"85", X"0c", X"81", X"d0", X"0c", 
    X"22", X"c0", X"0c", X"85", X"81", X"0c", X"ad", X"82", 
    X"ae", X"83", X"af", X"f0", X"74", X"24", X"2d", X"fa", 
    X"e4", X"3e", X"fb", X"8f", X"04", X"8a", X"82", X"8b", 
    X"83", X"8c", X"f0", X"12", X"70", X"5a", X"70", X"03", 
    X"02", X"44", X"2c", X"74", X"06", X"2d", X"fa", X"e4", 
    X"3e", X"fb", X"8f", X"04", X"74", X"03", X"2a", X"fa", 
    X"e4", X"3b", X"fb", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"12", X"70", X"5a", X"fa", X"a3", X"12", X"70", 
    X"5a", X"fb", X"a3", X"12", X"70", X"5a", X"fc", X"c0", 
    X"07", X"c0", X"06", X"c0", X"05", X"c0", X"04", X"c0", 
    X"03", X"c0", X"02", X"e5", X"0c", X"24", X"fb", X"f8", 
    X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"12", X"48", X"02", X"15", X"81", X"15", X"81", 
    X"15", X"81", X"d0", X"02", X"d0", X"03", X"d0", X"04", 
    X"d0", X"05", X"d0", X"06", X"d0", X"07", X"74", X"06", 
    X"2d", X"fd", X"e4", X"3e", X"fe", X"74", X"03", X"2d", 
    X"fd", X"e4", X"3e", X"fe", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"ea", X"12", X"66", X"a0", X"a3", X"eb", 
    X"12", X"66", X"a0", X"a3", X"ec", X"12", X"66", X"a0", 
    X"7f", X"01", X"80", X"02", X"7f", X"00", X"8f", X"82", 
    X"d0", X"0c", X"22", X"ad", X"82", X"ae", X"83", X"af", 
    X"f0", X"c0", X"e0", X"c0", X"a8", X"c2", X"af", X"74", 
    X"24", X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fd", 
    X"d0", X"e0", X"53", X"e0", X"80", X"e5", X"e0", X"42", 
    X"a8", X"d0", X"e0", X"8d", X"82", X"22", X"ad", X"82", 
    X"ae", X"83", X"af", X"f0", X"c0", X"e0", X"c0", X"a8", 
    X"c2", X"af", X"74", X"25", X"2d", X"fa", X"e4", X"3e", 
    X"fb", X"8f", X"04", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"12", X"70", X"5a", X"fa", X"74", X"24", X"2d", 
    X"fd", X"e4", X"3e", X"fe", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"70", X"5a", X"fd", X"ea", X"c3", 
    X"9d", X"fa", X"d0", X"e0", X"53", X"e0", X"80", X"e5", 
    X"e0", X"42", X"a8", X"d0", X"e0", X"8a", X"82", X"22", 
    X"ad", X"82", X"ae", X"83", X"af", X"f0", X"74", X"24", 
    X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"70", X"5a", X"f5", X"82", 
    X"22", X"12", X"62", X"2d", X"22", X"c0", X"0c", X"85", 
    X"81", X"0c", X"c0", X"82", X"c0", X"83", X"c0", X"f0", 
    X"e5", X"81", X"24", X"0a", X"f5", X"81", X"a8", X"0c", 
    X"08", X"74", X"24", X"26", X"fa", X"e4", X"08", X"36", 
    X"fb", X"08", X"86", X"04", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"e5", X"0c", X"24", X"0d", X"f8", X"12", 
    X"70", X"5a", X"f6", X"a8", X"0c", X"08", X"e5", X"0c", 
    X"24", X"04", X"f9", X"74", X"26", X"26", X"f7", X"e4", 
    X"08", X"36", X"09", X"f7", X"08", X"09", X"e6", X"f7", 
    X"e5", X"0c", X"24", X"04", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"fe", X"70", X"03", X"02", X"47", X"e9", X"e5", X"0c", 
    X"24", X"fa", X"f8", X"e6", X"60", X"03", X"02", X"46", 
    X"73", X"c0", X"02", X"c0", X"03", X"c0", X"04", X"8e", 
    X"04", X"7d", X"00", X"a8", X"0c", X"08", X"e5", X"0c", 
    X"24", X"07", X"f9", X"74", X"03", X"26", X"f7", X"e4", 
    X"08", X"36", X"09", X"f7", X"08", X"09", X"e6", X"f7", 
    X"e5", X"0c", X"24", X"07", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"fa", X"a3", X"12", X"70", X"5a", X"fb", X"a3", X"12", 
    X"70", X"5a", X"ff", X"c0", X"04", X"c0", X"03", X"c0", 
    X"02", X"c0", X"04", X"c0", X"05", X"e5", X"0c", X"24", 
    X"fb", X"f8", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"08", X"e6", X"c0", X"e0", X"8a", X"82", X"8b", 
    X"83", X"8f", X"f0", X"12", X"67", X"03", X"e5", X"81", 
    X"24", X"fb", X"f5", X"81", X"d0", X"02", X"d0", X"03", 
    X"d0", X"04", X"e5", X"0c", X"24", X"07", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"12", 
    X"70", X"5a", X"fc", X"a3", X"12", X"70", X"5a", X"fd", 
    X"a3", X"12", X"70", X"5a", X"ff", X"e5", X"0c", X"24", 
    X"04", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"12", X"70", X"5a", X"fb", X"e5", X"0c", 
    X"24", X"0a", X"f8", X"eb", X"2c", X"f6", X"e4", X"3d", 
    X"08", X"f6", X"08", X"a6", X"07", X"e5", X"0c", X"24", 
    X"07", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"e5", X"0c", X"24", X"0a", X"f9", X"e7", 
    X"12", X"66", X"a0", X"a3", X"09", X"e7", X"12", X"66", 
    X"a0", X"a3", X"09", X"e7", X"12", X"66", X"a0", X"a8", 
    X"0c", X"08", X"74", X"06", X"26", X"fa", X"e4", X"08", 
    X"36", X"fb", X"08", X"86", X"07", X"8a", X"82", X"8b", 
    X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fa", X"a3", 
    X"12", X"70", X"5a", X"fb", X"a3", X"12", X"70", X"5a", 
    X"ff", X"e5", X"0c", X"24", X"0a", X"f8", X"c0", X"02", 
    X"c0", X"03", X"c0", X"07", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"00", X"11", X"15", 
    X"81", X"15", X"81", X"15", X"81", X"d0", X"04", X"d0", 
    X"03", X"d0", X"02", X"50", X"03", X"02", X"47", X"e9", 
    X"c0", X"02", X"c0", X"03", X"c0", X"04", X"a8", X"0c", 
    X"08", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"70", X"5a", X"fc", X"a3", X"12", X"70", 
    X"5a", X"fd", X"a3", X"12", X"70", X"5a", X"ff", X"e5", 
    X"0c", X"24", X"07", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"ec", X"12", X"66", X"a0", 
    X"a3", X"ed", X"12", X"66", X"a0", X"a3", X"ef", X"12", 
    X"66", X"a0", X"d0", X"04", X"d0", X"03", X"d0", X"02", 
    X"02", X"47", X"e9", X"c0", X"02", X"c0", X"03", X"c0", 
    X"04", X"7f", X"00", X"a8", X"0c", X"08", X"e5", X"0c", 
    X"24", X"0a", X"f9", X"74", X"06", X"26", X"f7", X"e4", 
    X"08", X"36", X"09", X"f7", X"08", X"09", X"e6", X"f7", 
    X"e5", X"0c", X"24", X"0a", X"f8", X"e5", X"0c", X"24", 
    X"07", X"f9", X"74", X"03", X"26", X"f7", X"e4", X"08", 
    X"36", X"09", X"f7", X"08", X"09", X"e6", X"f7", X"e5", 
    X"0c", X"24", X"07", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", X"fb", 
    X"a3", X"12", X"70", X"5a", X"fc", X"a3", X"12", X"70", 
    X"5a", X"fd", X"c0", X"04", X"c0", X"03", X"c0", X"02", 
    X"c0", X"06", X"c0", X"07", X"e5", X"0c", X"24", X"fb", 
    X"f8", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", 
    X"08", X"e6", X"c0", X"e0", X"8b", X"82", X"8c", X"83", 
    X"8d", X"f0", X"12", X"67", X"03", X"e5", X"81", X"24", 
    X"fb", X"f5", X"81", X"d0", X"02", X"d0", X"03", X"d0", 
    X"04", X"e5", X"0c", X"24", X"07", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"70", 
    X"5a", X"fd", X"a3", X"12", X"70", X"5a", X"fe", X"a3", 
    X"12", X"70", X"5a", X"ff", X"e5", X"0c", X"24", X"04", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"70", X"5a", X"fc", X"7b", X"00", X"ed", 
    X"c3", X"9c", X"fd", X"ee", X"9b", X"fe", X"e5", X"0c", 
    X"24", X"07", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"ed", X"12", X"66", X"a0", X"a3", 
    X"ee", X"12", X"66", X"a0", X"a3", X"ef", X"12", X"66", 
    X"a0", X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", X"fa", 
    X"a3", X"12", X"70", X"5a", X"fb", X"a3", X"12", X"70", 
    X"5a", X"fc", X"c0", X"02", X"c0", X"03", X"c0", X"04", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"00", 
    X"11", X"15", X"81", X"15", X"81", X"15", X"81", X"d0", 
    X"04", X"d0", X"03", X"d0", X"02", X"50", X"5c", X"c0", 
    X"02", X"c0", X"03", X"c0", X"04", X"e5", X"0c", X"24", 
    X"0a", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"12", X"70", X"5a", X"fd", X"a3", X"12", 
    X"70", X"5a", X"fe", X"a3", X"12", X"70", X"5a", X"ff", 
    X"e5", X"0c", X"24", X"04", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"fc", X"7b", X"00", X"ed", X"c3", X"9c", X"fd", X"ee", 
    X"9b", X"fe", X"e5", X"0c", X"24", X"07", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"ed", 
    X"12", X"66", X"a0", X"a3", X"ee", X"12", X"66", X"a0", 
    X"a3", X"ef", X"12", X"66", X"a0", X"d0", X"04", X"d0", 
    X"03", X"d0", X"02", X"e5", X"0c", X"24", X"fa", X"f8", 
    X"b6", X"02", X"0e", X"e5", X"0c", X"24", X"0d", X"f8", 
    X"e6", X"60", X"06", X"e5", X"0c", X"24", X"0d", X"f8", 
    X"16", X"e5", X"0c", X"24", X"0d", X"f8", X"e6", X"04", 
    X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"12", X"66", 
    X"a0", X"75", X"82", X"00", X"85", X"0c", X"81", X"d0", 
    X"0c", X"22", X"c0", X"0c", X"85", X"81", X"0c", X"c0", 
    X"82", X"c0", X"83", X"c0", X"f0", X"e5", X"81", X"24", 
    X"04", X"f5", X"81", X"a8", X"0c", X"08", X"74", X"26", 
    X"26", X"fa", X"e4", X"08", X"36", X"fb", X"08", X"86", 
    X"04", X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"e5", 
    X"0c", X"24", X"04", X"f8", X"12", X"70", X"5a", X"f6", 
    X"e5", X"0c", X"24", X"04", X"f8", X"e6", X"70", X"03", 
    X"02", X"49", X"4c", X"c0", X"02", X"c0", X"03", X"c0", 
    X"04", X"a8", X"0c", X"08", X"74", X"06", X"26", X"fa", 
    X"e4", X"08", X"36", X"fb", X"08", X"86", X"04", X"e5", 
    X"0c", X"24", X"05", X"f8", X"74", X"03", X"2a", X"f6", 
    X"e4", X"3b", X"08", X"f6", X"08", X"a6", X"04", X"e5", 
    X"0c", X"24", X"05", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", X"fd", 
    X"a3", X"12", X"70", X"5a", X"fe", X"a3", X"12", X"70", 
    X"5a", X"ff", X"e5", X"0c", X"24", X"04", X"f8", X"e6", 
    X"2d", X"fd", X"e4", X"3e", X"fe", X"e5", X"0c", X"24", 
    X"05", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"ed", X"12", X"66", X"a0", X"a3", X"ee", 
    X"12", X"66", X"a0", X"a3", X"ef", X"12", X"66", X"a0", 
    X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"12", X"70", 
    X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"fb", X"a3", 
    X"12", X"70", X"5a", X"fc", X"c0", X"02", X"c0", X"03", 
    X"c0", X"04", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"00", X"11", X"15", X"81", X"15", X"81", X"15", 
    X"81", X"d0", X"04", X"d0", X"03", X"d0", X"02", X"40", 
    X"34", X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", X"fd", 
    X"a3", X"12", X"70", X"5a", X"fe", X"a3", X"12", X"70", 
    X"5a", X"ff", X"e5", X"0c", X"24", X"05", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"ed", 
    X"12", X"66", X"a0", X"a3", X"ee", X"12", X"66", X"a0", 
    X"a3", X"ef", X"12", X"66", X"a0", X"8a", X"82", X"8b", 
    X"83", X"8c", X"f0", X"12", X"70", X"5a", X"fa", X"7f", 
    X"00", X"e5", X"0c", X"24", X"05", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"70", 
    X"5a", X"fc", X"a3", X"12", X"70", X"5a", X"fd", X"a3", 
    X"12", X"70", X"5a", X"fe", X"c0", X"02", X"c0", X"07", 
    X"c0", X"04", X"c0", X"05", X"c0", X"06", X"e5", X"0c", 
    X"24", X"fb", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"67", X"03", X"e5", X"81", 
    X"24", X"fb", X"f5", X"81", X"85", X"0c", X"81", X"d0", 
    X"0c", X"22", X"c0", X"0c", X"85", X"81", X"0c", X"c0", 
    X"82", X"c0", X"83", X"c0", X"f0", X"e5", X"81", X"24", 
    X"04", X"f5", X"81", X"c0", X"e0", X"c0", X"a8", X"c2", 
    X"af", X"a8", X"0c", X"08", X"74", X"28", X"26", X"fa", 
    X"e4", X"08", X"36", X"fb", X"08", X"86", X"04", X"8a", 
    X"82", X"8b", X"83", X"8c", X"f0", X"e5", X"0c", X"24", 
    X"07", X"f8", X"12", X"70", X"5a", X"f6", X"a8", X"0c", 
    X"08", X"e5", X"0c", X"24", X"04", X"f9", X"74", X"18", 
    X"26", X"f7", X"e4", X"08", X"36", X"09", X"f7", X"08", 
    X"09", X"e6", X"f7", X"e5", X"0c", X"24", X"07", X"f8", 
    X"c3", X"74", X"80", X"86", X"f0", X"63", X"f0", X"80", 
    X"95", X"f0", X"50", X"50", X"e5", X"0c", X"24", X"04", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"70", X"5a", X"60", X"3e", X"a8", X"0c", 
    X"08", X"74", X"18", X"26", X"fd", X"e4", X"08", X"36", 
    X"fe", X"08", X"86", X"07", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"c0", X"04", X"c0", X"03", X"c0", X"02", 
    X"12", X"10", X"57", X"e5", X"82", X"d0", X"02", X"d0", 
    X"03", X"d0", X"04", X"60", X"0f", X"c0", X"04", X"c0", 
    X"03", X"c0", X"02", X"12", X"14", X"4d", X"d0", X"02", 
    X"d0", X"03", X"d0", X"04", X"e5", X"0c", X"24", X"07", 
    X"f8", X"16", X"80", X"9f", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"74", X"ff", X"12", X"66", X"a0", X"d0", 
    X"e0", X"53", X"e0", X"80", X"e5", X"e0", X"42", X"a8", 
    X"d0", X"e0", X"c0", X"e0", X"c0", X"a8", X"c2", X"af", 
    X"a8", X"0c", X"08", X"74", X"27", X"26", X"fd", X"e4", 
    X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fc", 
    X"a8", X"0c", X"08", X"e5", X"0c", X"24", X"04", X"f9", 
    X"74", X"0c", X"26", X"f7", X"e4", X"08", X"36", X"09", 
    X"f7", X"08", X"09", X"e6", X"f7", X"c3", X"74", X"80", 
    X"8c", X"f0", X"63", X"f0", X"80", X"95", X"f0", X"50", 
    X"5f", X"e5", X"0c", X"24", X"04", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"70", 
    X"5a", X"60", X"4d", X"c0", X"05", X"c0", X"06", X"c0", 
    X"07", X"a8", X"0c", X"08", X"74", X"0c", X"26", X"fa", 
    X"e4", X"08", X"36", X"fb", X"08", X"86", X"07", X"8a", 
    X"82", X"8b", X"83", X"8f", X"f0", X"c0", X"07", X"c0", 
    X"06", X"c0", X"05", X"c0", X"04", X"12", X"10", X"57", 
    X"e5", X"82", X"d0", X"04", X"d0", X"05", X"d0", X"06", 
    X"d0", X"07", X"d0", X"07", X"d0", X"06", X"d0", X"05", 
    X"60", X"13", X"c0", X"07", X"c0", X"06", X"c0", X"05", 
    X"c0", X"04", X"12", X"14", X"4d", X"d0", X"04", X"d0", 
    X"05", X"d0", X"06", X"d0", X"07", X"1c", X"80", X"95", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"74", X"ff", 
    X"12", X"66", X"a0", X"d0", X"e0", X"53", X"e0", X"80", 
    X"e5", X"e0", X"42", X"a8", X"d0", X"e0", X"85", X"0c", 
    X"81", X"d0", X"0c", X"22", X"ad", X"82", X"ae", X"83", 
    X"af", X"f0", X"c0", X"e0", X"c0", X"a8", X"c2", X"af", 
    X"74", X"24", X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"70", X"04", X"7f", X"01", X"80", X"02", X"7f", X"00", 
    X"d0", X"e0", X"53", X"e0", X"80", X"e5", X"e0", X"42", 
    X"a8", X"d0", X"e0", X"8f", X"82", X"22", X"ad", X"82", 
    X"ae", X"83", X"af", X"f0", X"74", X"24", X"2d", X"fd", 
    X"e4", X"3e", X"fe", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"12", X"70", X"5a", X"70", X"04", X"7f", X"01", 
    X"80", X"02", X"7f", X"00", X"8f", X"82", X"22", X"ad", 
    X"82", X"ae", X"83", X"af", X"f0", X"c0", X"e0", X"c0", 
    X"a8", X"c2", X"af", X"74", X"24", X"2d", X"fa", X"e4", 
    X"3e", X"fb", X"8f", X"04", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"12", X"70", X"5a", X"fa", X"74", X"25", 
    X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fd", X"ea", 
    X"b5", X"05", X"04", X"7f", X"01", X"80", X"02", X"7f", 
    X"00", X"d0", X"e0", X"53", X"e0", X"80", X"e5", X"e0", 
    X"42", X"a8", X"d0", X"e0", X"8f", X"82", X"22", X"ad", 
    X"82", X"ae", X"83", X"af", X"f0", X"74", X"24", X"2d", 
    X"fa", X"e4", X"3e", X"fb", X"8f", X"04", X"8a", X"82", 
    X"8b", X"83", X"8c", X"f0", X"12", X"70", X"5a", X"fa", 
    X"74", X"25", X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"fd", X"ea", X"b5", X"05", X"04", X"7f", X"01", X"80", 
    X"02", X"7f", X"00", X"8f", X"82", X"22", X"c0", X"0c", 
    X"e5", X"81", X"f5", X"0c", X"24", X"06", X"f5", X"81", 
    X"ae", X"82", X"af", X"83", X"e5", X"0c", X"24", X"fb", 
    X"f8", X"b6", X"01", X"09", X"e5", X"0c", X"24", X"06", 
    X"f8", X"76", X"01", X"80", X"07", X"e5", X"0c", X"24", 
    X"06", X"f8", X"76", X"00", X"e5", X"0c", X"24", X"fc", 
    X"f8", X"e6", X"08", X"46", X"70", X"0a", X"e5", X"0c", 
    X"24", X"fc", X"f8", X"76", X"01", X"08", X"76", X"00", 
    X"a8", X"0c", X"08", X"74", X"01", X"2e", X"f6", X"e4", 
    X"3f", X"08", X"f6", X"a8", X"0c", X"08", X"74", X"12", 
    X"26", X"fb", X"e4", X"08", X"36", X"fc", X"8b", X"82", 
    X"8c", X"83", X"12", X"61", X"84", X"aa", X"82", X"ab", 
    X"83", X"ac", X"f0", X"e5", X"0c", X"24", X"03", X"f8", 
    X"a6", X"02", X"08", X"a6", X"03", X"08", X"a6", X"04", 
    X"e5", X"0c", X"24", X"03", X"f8", X"e6", X"08", X"46", 
    X"60", X"50", X"e5", X"0c", X"24", X"03", X"f8", X"74", 
    X"12", X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", 
    X"86", X"07", X"e5", X"0c", X"24", X"03", X"f8", X"86", 
    X"02", X"08", X"86", X"03", X"08", X"86", X"04", X"e5", 
    X"0c", X"24", X"06", X"f8", X"e6", X"c0", X"e0", X"e5", 
    X"0c", X"24", X"fc", X"f8", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"a8", X"0c", X"08", X"e6", X"c0", 
    X"e0", X"08", X"e6", X"c0", X"e0", X"c0", X"05", X"c0", 
    X"06", X"c0", X"07", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"12", X"60", X"d6", X"e5", X"81", X"24", X"f8", 
    X"f5", X"81", X"e5", X"0c", X"24", X"03", X"f8", X"86", 
    X"02", X"08", X"86", X"03", X"08", X"86", X"04", X"8a", 
    X"82", X"8b", X"83", X"8c", X"f0", X"85", X"0c", X"81", 
    X"d0", X"0c", X"22", X"ad", X"82", X"ae", X"83", X"af", 
    X"f0", X"8d", X"02", X"8e", X"03", X"8f", X"04", X"74", 
    X"11", X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"20", 
    X"e1", X"11", X"8a", X"05", X"8b", X"06", X"8c", X"07", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"62", 
    X"2d", X"80", X"18", X"74", X"12", X"c0", X"e0", X"e4", 
    X"c0", X"e0", X"c0", X"e0", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"12", X"66", X"db", X"15", X"81", X"15", 
    X"81", X"15", X"81", X"22", X"c0", X"0c", X"85", X"81", 
    X"0c", X"c0", X"82", X"c0", X"83", X"c0", X"f0", X"05", 
    X"81", X"05", X"81", X"05", X"81", X"7f", X"00", X"c0", 
    X"e0", X"c0", X"a8", X"c2", X"af", X"a8", X"0c", X"08", 
    X"74", X"08", X"26", X"fa", X"e4", X"08", X"36", X"fb", 
    X"08", X"86", X"04", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"12", X"70", X"5a", X"fa", X"a3", X"12", X"70", 
    X"5a", X"fb", X"a3", X"12", X"70", X"5a", X"fc", X"ea", 
    X"4b", X"60", X"03", X"02", X"4d", X"e2", X"a8", X"0c", 
    X"08", X"74", X"0b", X"26", X"fa", X"e4", X"08", X"36", 
    X"fb", X"08", X"86", X"04", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"12", X"70", X"5a", X"fa", X"a3", X"12", 
    X"70", X"5a", X"fb", X"a3", X"12", X"70", X"5a", X"fc", 
    X"ea", X"4b", X"60", X"03", X"02", X"4d", X"e2", X"a8", 
    X"0c", X"08", X"74", X"11", X"26", X"fa", X"e4", X"08", 
    X"36", X"fb", X"08", X"86", X"04", X"8a", X"82", X"8b", 
    X"83", X"8c", X"f0", X"e5", X"0c", X"24", X"04", X"f8", 
    X"12", X"70", X"5a", X"f6", X"a8", X"0c", X"08", X"74", 
    X"06", X"26", X"fb", X"e4", X"08", X"36", X"fc", X"08", 
    X"86", X"07", X"8b", X"82", X"8c", X"83", X"8f", X"f0", 
    X"12", X"70", X"5a", X"fb", X"a3", X"12", X"70", X"5a", 
    X"fc", X"a8", X"0c", X"08", X"74", X"04", X"26", X"fd", 
    X"e4", X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"e5", X"0c", X"24", 
    X"05", X"f8", X"12", X"70", X"5a", X"f6", X"a3", X"12", 
    X"70", X"5a", X"08", X"f6", X"a8", X"0c", X"08", X"74", 
    X"0e", X"26", X"fa", X"e4", X"08", X"36", X"fe", X"08", 
    X"86", X"07", X"8a", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"70", X"5a", X"fa", X"a3", X"12", X"70", X"5a", 
    X"fe", X"a3", X"12", X"70", X"5a", X"ff", X"e5", X"0c", 
    X"24", X"04", X"f8", X"e6", X"c0", X"e0", X"c0", X"03", 
    X"c0", X"04", X"e5", X"0c", X"24", X"05", X"f8", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"c0", X"02", 
    X"c0", X"06", X"c0", X"07", X"a8", X"0c", X"08", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"12", 
    X"60", X"d6", X"e5", X"81", X"24", X"f8", X"f5", X"81", 
    X"7f", X"01", X"d0", X"e0", X"53", X"e0", X"80", X"e5", 
    X"e0", X"42", X"a8", X"d0", X"e0", X"8f", X"82", X"85", 
    X"0c", X"81", X"d0", X"0c", X"22", X"c0", X"0c", X"85", 
    X"81", X"0c", X"ad", X"82", X"ae", X"83", X"af", X"f0", 
    X"e5", X"0c", X"24", X"fc", X"f8", X"e6", X"08", X"46", 
    X"70", X"0a", X"e5", X"0c", X"24", X"fc", X"f8", X"76", 
    X"01", X"08", X"76", X"00", X"74", X"04", X"2d", X"fa", 
    X"e4", X"3e", X"fb", X"8f", X"04", X"8a", X"82", X"8b", 
    X"83", X"8c", X"f0", X"12", X"70", X"5a", X"fa", X"a3", 
    X"12", X"70", X"5a", X"fb", X"e5", X"0c", X"24", X"fc", 
    X"f8", X"c3", X"ea", X"96", X"eb", X"08", X"96", X"40", 
    X"20", X"74", X"06", X"2d", X"fd", X"e4", X"3e", X"fe", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"e5", X"0c", 
    X"24", X"fc", X"f8", X"e6", X"12", X"66", X"a0", X"a3", 
    X"08", X"e6", X"12", X"66", X"a0", X"7f", X"01", X"80", 
    X"02", X"7f", X"00", X"8f", X"82", X"d0", X"0c", X"22", 
    X"c0", X"0c", X"85", X"81", X"0c", X"c0", X"82", X"c0", 
    X"83", X"c0", X"f0", X"05", X"81", X"05", X"81", X"a8", 
    X"0c", X"08", X"74", X"04", X"26", X"fb", X"e4", X"08", 
    X"36", X"fa", X"08", X"86", X"04", X"8b", X"82", X"8a", 
    X"83", X"8c", X"f0", X"12", X"70", X"5a", X"fb", X"a3", 
    X"12", X"70", X"5a", X"fc", X"a8", X"0c", X"08", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"12", 
    X"70", X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"ff", 
    X"e5", X"0c", X"24", X"04", X"f8", X"ea", X"2b", X"f6", 
    X"ef", X"3c", X"08", X"f6", X"a8", X"0c", X"08", X"74", 
    X"02", X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", 
    X"86", X"07", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"70", X"5a", X"fd", X"a3", X"12", X"70", X"5a", 
    X"fe", X"e5", X"0c", X"24", X"04", X"f8", X"e6", X"c3", 
    X"9d", X"fd", X"08", X"e6", X"9e", X"fe", X"ed", X"24", 
    X"ff", X"ff", X"ee", X"34", X"ff", X"fe", X"c3", X"ef", 
    X"9b", X"ee", X"9c", X"40", X"07", X"ef", X"c3", X"9b", 
    X"ff", X"ee", X"9c", X"fe", X"8f", X"82", X"8e", X"83", 
    X"85", X"0c", X"81", X"d0", X"0c", X"22", X"12", X"60", 
    X"56", X"22", X"c0", X"0c", X"e5", X"81", X"f5", X"0c", 
    X"24", X"0d", X"f5", X"81", X"ad", X"82", X"ae", X"83", 
    X"af", X"f0", X"e5", X"0c", X"24", X"04", X"f8", X"a6", 
    X"05", X"08", X"a6", X"06", X"08", X"a6", X"07", X"e5", 
    X"0c", X"24", X"07", X"f8", X"e4", X"f6", X"08", X"f6", 
    X"e5", X"0c", X"24", X"f9", X"f8", X"e5", X"0c", X"24", 
    X"09", X"f9", X"e6", X"f7", X"08", X"09", X"e6", X"f7", 
    X"74", X"11", X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"fd", X"30", X"e0", X"0d", X"e5", X"0c", X"24", X"09", 
    X"f8", X"74", X"02", X"26", X"f6", X"e4", X"08", X"36", 
    X"f6", X"e5", X"0c", X"24", X"f7", X"f8", X"e6", X"08", 
    X"46", X"70", X"03", X"02", X"50", X"8d", X"e5", X"0c", 
    X"24", X"0b", X"ff", X"fc", X"7d", X"00", X"7e", X"40", 
    X"8c", X"82", X"8d", X"83", X"8e", X"f0", X"c0", X"07", 
    X"12", X"12", X"dd", X"d0", X"07", X"a8", X"0c", X"08", 
    X"a6", X"07", X"c0", X"e0", X"c0", X"a8", X"c2", X"af", 
    X"e5", X"0c", X"24", X"04", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"4e", X"60", 
    X"ae", X"82", X"af", X"83", X"e5", X"0c", X"24", X"07", 
    X"f8", X"a6", X"06", X"08", X"a6", X"07", X"e5", X"0c", 
    X"24", X"07", X"f8", X"e5", X"0c", X"24", X"09", X"f9", 
    X"c3", X"e6", X"97", X"08", X"e6", X"09", X"97", X"50", 
    X"44", X"90", X"00", X"00", X"75", X"f0", X"00", X"12", 
    X"21", X"e1", X"e5", X"0c", X"24", X"04", X"f8", X"74", 
    X"0b", X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", 
    X"86", X"07", X"c0", X"07", X"c0", X"06", X"c0", X"05", 
    X"12", X"15", X"47", X"aa", X"82", X"ab", X"83", X"ac", 
    X"f0", X"d0", X"05", X"d0", X"06", X"d0", X"07", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"ea", X"12", X"66", 
    X"a0", X"a3", X"eb", X"12", X"66", X"a0", X"a3", X"ec", 
    X"12", X"66", X"a0", X"80", X"0e", X"d0", X"e0", X"53", 
    X"e0", X"80", X"e5", X"e0", X"42", X"a8", X"d0", X"e0", 
    X"02", X"50", X"8d", X"d0", X"e0", X"53", X"e0", X"80", 
    X"e5", X"e0", X"42", X"a8", X"d0", X"e0", X"c0", X"07", 
    X"c0", X"06", X"c0", X"05", X"e5", X"0c", X"24", X"f7", 
    X"f8", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", 
    X"e4", X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", 
    X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", X"90", 
    X"00", X"00", X"e4", X"f5", X"f0", X"12", X"17", X"6d", 
    X"e5", X"81", X"24", X"f7", X"f5", X"81", X"d0", X"05", 
    X"d0", X"06", X"d0", X"07", X"7a", X"00", X"7b", X"00", 
    X"7c", X"00", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"ea", X"12", X"66", X"a0", X"a3", X"eb", X"12", X"66", 
    X"a0", X"a3", X"ec", X"12", X"66", X"a0", X"e5", X"0c", 
    X"24", X"f7", X"ff", X"7e", X"00", X"7d", X"40", X"a8", 
    X"0c", X"08", X"86", X"02", X"7b", X"00", X"7c", X"40", 
    X"c0", X"07", X"c0", X"06", X"c0", X"05", X"8a", X"82", 
    X"8b", X"83", X"8c", X"f0", X"12", X"13", X"4e", X"af", 
    X"82", X"15", X"81", X"15", X"81", X"15", X"81", X"ef", 
    X"70", X"03", X"02", X"4f", X"7a", X"e5", X"0c", X"24", 
    X"07", X"f8", X"e6", X"08", X"46", X"70", X"1e", X"e5", 
    X"0c", X"24", X"04", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"4e", X"60", X"ae", 
    X"82", X"af", X"83", X"e5", X"0c", X"24", X"07", X"f8", 
    X"a6", X"06", X"08", X"a6", X"07", X"e5", X"0c", X"24", 
    X"09", X"f8", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"e5", X"0c", X"24", X"07", X"f8", X"e6", X"c0", 
    X"e0", X"08", X"e6", X"c0", X"e0", X"e5", X"0c", X"24", 
    X"f9", X"f8", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"e5", X"0c", X"24", X"fb", X"f8", X"e6", X"c0", 
    X"e0", X"08", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"e5", X"0c", X"24", X"04", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"53", 
    X"65", X"ae", X"82", X"af", X"83", X"e5", X"81", X"24", 
    X"f7", X"f5", X"81", X"a8", X"0c", X"08", X"08", X"a6", 
    X"06", X"08", X"a6", X"07", X"ee", X"4f", X"70", X"03", 
    X"02", X"51", X"d7", X"e5", X"0c", X"24", X"04", X"f8", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"12", X"60", X"56", X"ae", X"82", X"af", X"83", X"e5", 
    X"0c", X"24", X"04", X"f8", X"74", X"06", X"26", X"fb", 
    X"e4", X"08", X"36", X"fc", X"08", X"86", X"05", X"8b", 
    X"82", X"8c", X"83", X"8d", X"f0", X"12", X"70", X"5a", 
    X"fb", X"a3", X"12", X"70", X"5a", X"fc", X"c3", X"ee", 
    X"9b", X"ef", X"9c", X"50", X"03", X"02", X"51", X"d7", 
    X"12", X"09", X"4a", X"e5", X"0c", X"24", X"04", X"f8", 
    X"74", X"08", X"26", X"fb", X"e4", X"08", X"36", X"fc", 
    X"08", X"86", X"06", X"8b", X"82", X"8c", X"83", X"8e", 
    X"f0", X"12", X"70", X"5a", X"fa", X"a3", X"12", X"70", 
    X"5a", X"fd", X"a3", X"12", X"70", X"5a", X"ea", X"4d", 
    X"60", X"5a", X"8b", X"82", X"8c", X"83", X"8e", X"f0", 
    X"12", X"70", X"5a", X"fa", X"a3", X"12", X"70", X"5a", 
    X"fd", X"a3", X"12", X"70", X"5a", X"ff", X"c0", X"06", 
    X"c0", X"04", X"c0", X"03", X"e4", X"c0", X"e0", X"c0", 
    X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", 
    X"e0", X"c0", X"e0", X"c0", X"e0", X"8a", X"82", X"8d", 
    X"83", X"8f", X"f0", X"12", X"19", X"e0", X"e5", X"81", 
    X"24", X"f8", X"f5", X"81", X"d0", X"03", X"d0", X"04", 
    X"d0", X"06", X"7a", X"00", X"7d", X"00", X"7f", X"00", 
    X"8b", X"82", X"8c", X"83", X"8e", X"f0", X"ea", X"12", 
    X"66", X"a0", X"a3", X"ed", X"12", X"66", X"a0", X"a3", 
    X"ef", X"12", X"66", X"a0", X"12", X"09", X"52", X"a8", 
    X"0c", X"08", X"08", X"86", X"82", X"08", X"86", X"83", 
    X"85", X"0c", X"81", X"d0", X"0c", X"22", X"c0", X"0c", 
    X"e5", X"81", X"f5", X"0c", X"24", X"05", X"f5", X"81", 
    X"ad", X"82", X"ae", X"83", X"af", X"f0", X"e5", X"0c", 
    X"24", X"03", X"f8", X"a6", X"05", X"08", X"a6", X"06", 
    X"08", X"a6", X"07", X"e5", X"0c", X"24", X"f9", X"f8", 
    X"86", X"04", X"08", X"86", X"03", X"74", X"11", X"2d", 
    X"fd", X"e4", X"3e", X"fe", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"70", X"5a", X"30", X"e0", X"07", 
    X"74", X"02", X"2c", X"fc", X"e4", X"3b", X"fb", X"e5", 
    X"0c", X"24", X"03", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"c0", X"04", X"c0", X"03", 
    X"12", X"4e", X"60", X"ae", X"82", X"af", X"83", X"c0", 
    X"06", X"c0", X"07", X"e5", X"0c", X"24", X"f9", X"f8", 
    X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"e5", 
    X"0c", X"24", X"fb", X"f8", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"e5", 
    X"0c", X"24", X"03", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"53", X"65", X"ae", 
    X"82", X"af", X"83", X"e5", X"81", X"24", X"f7", X"f5", 
    X"81", X"a8", X"0c", X"08", X"a6", X"06", X"08", X"a6", 
    X"07", X"ee", X"4f", X"70", X"03", X"02", X"53", X"57", 
    X"e5", X"0c", X"24", X"03", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"60", X"56", 
    X"ae", X"82", X"af", X"83", X"e5", X"0c", X"24", X"03", 
    X"f8", X"74", X"06", X"26", X"fb", X"e4", X"08", X"36", 
    X"fc", X"08", X"86", X"05", X"8b", X"82", X"8c", X"83", 
    X"8d", X"f0", X"12", X"70", X"5a", X"fb", X"a3", X"12", 
    X"70", X"5a", X"fc", X"c3", X"ee", X"9b", X"ef", X"9c", 
    X"50", X"03", X"02", X"53", X"57", X"e5", X"0c", X"24", 
    X"03", X"f8", X"74", X"08", X"26", X"fb", X"e4", X"08", 
    X"36", X"fc", X"08", X"86", X"06", X"8b", X"82", X"8c", 
    X"83", X"8e", X"f0", X"12", X"70", X"5a", X"fa", X"a3", 
    X"12", X"70", X"5a", X"fd", X"a3", X"12", X"70", X"5a", 
    X"ff", X"ea", X"4d", X"60", X"6a", X"8b", X"82", X"8c", 
    X"83", X"8e", X"f0", X"12", X"70", X"5a", X"fa", X"a3", 
    X"12", X"70", X"5a", X"fd", X"a3", X"12", X"70", X"5a", 
    X"ff", X"c0", X"06", X"c0", X"04", X"c0", X"03", X"e5", 
    X"0c", X"24", X"f6", X"f8", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"e4", 
    X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", 
    X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", 
    X"8a", X"82", X"8d", X"83", X"8f", X"f0", X"12", X"1c", 
    X"d7", X"e5", X"81", X"24", X"f5", X"f5", X"81", X"d0", 
    X"03", X"d0", X"04", X"d0", X"06", X"7a", X"00", X"7d", 
    X"00", X"7f", X"00", X"8b", X"82", X"8c", X"83", X"8e", 
    X"f0", X"ea", X"12", X"66", X"a0", X"a3", X"ed", X"12", 
    X"66", X"a0", X"a3", X"ef", X"12", X"66", X"a0", X"a8", 
    X"0c", X"08", X"86", X"82", X"08", X"86", X"83", X"85", 
    X"0c", X"81", X"d0", X"0c", X"22", X"c0", X"0c", X"85", 
    X"81", X"0c", X"c0", X"82", X"c0", X"83", X"c0", X"f0", 
    X"e5", X"0c", X"24", X"f7", X"f8", X"e6", X"08", X"46", 
    X"70", X"04", X"fc", X"02", X"54", X"17", X"a8", X"0c", 
    X"08", X"74", X"11", X"26", X"fa", X"e4", X"08", X"36", 
    X"fb", X"08", X"86", X"07", X"8a", X"82", X"8b", X"83", 
    X"8f", X"f0", X"12", X"70", X"5a", X"fa", X"20", X"e0", 
    X"37", X"7c", X"01", X"e5", X"0c", X"24", X"f9", X"f8", 
    X"e5", X"0c", X"24", X"f7", X"f9", X"c3", X"e6", X"97", 
    X"08", X"e6", X"09", X"97", X"50", X"0c", X"e5", X"0c", 
    X"24", X"f9", X"f8", X"86", X"06", X"08", X"86", X"07", 
    X"80", X"0a", X"e5", X"0c", X"24", X"f7", X"f8", X"86", 
    X"06", X"08", X"86", X"07", X"e5", X"0c", X"24", X"f9", 
    X"f8", X"a6", X"06", X"08", X"a6", X"07", X"80", X"47", 
    X"e5", X"0c", X"24", X"f7", X"f8", X"e5", X"0c", X"24", 
    X"f5", X"f9", X"c3", X"e6", X"97", X"08", X"e6", X"09", 
    X"97", X"40", X"32", X"7c", X"01", X"e5", X"0c", X"24", 
    X"f9", X"ff", X"7e", X"00", X"7d", X"40", X"c0", X"04", 
    X"74", X"02", X"c0", X"e0", X"e4", X"c0", X"e0", X"c0", 
    X"07", X"c0", X"06", X"c0", X"05", X"a8", X"0c", X"08", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"12", X"5b", X"f4", X"e5", X"81", X"24", X"fb", X"f5", 
    X"81", X"d0", X"04", X"80", X"02", X"7c", X"00", X"ec", 
    X"60", X"39", X"e5", X"0c", X"24", X"fb", X"f8", X"86", 
    X"05", X"08", X"86", X"06", X"08", X"86", X"07", X"e5", 
    X"0c", X"24", X"f9", X"f8", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"c0", X"05", X"c0", X"06", X"c0", 
    X"07", X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"5b", X"f4", X"ae", 
    X"82", X"af", X"83", X"e5", X"81", X"24", X"fb", X"f5", 
    X"81", X"80", X"04", X"7e", X"00", X"7f", X"00", X"8e", 
    X"82", X"8f", X"83", X"85", X"0c", X"81", X"d0", X"0c", 
    X"22", X"c0", X"0c", X"e5", X"81", X"f5", X"0c", X"24", 
    X"09", X"f5", X"81", X"af", X"82", X"ae", X"83", X"ad", 
    X"f0", X"e5", X"0c", X"24", X"03", X"f8", X"a6", X"07", 
    X"08", X"a6", X"06", X"08", X"a6", X"05", X"a8", X"0c", 
    X"08", X"e4", X"f6", X"08", X"f6", X"74", X"11", X"2f", 
    X"fb", X"e4", X"3e", X"fc", X"8b", X"82", X"8c", X"83", 
    X"8d", X"f0", X"12", X"70", X"5a", X"fb", X"30", X"e0", 
    X"0c", X"e5", X"0c", X"24", X"08", X"f8", X"76", X"02", 
    X"08", X"76", X"00", X"80", X"09", X"e5", X"0c", X"24", 
    X"08", X"f8", X"e4", X"f6", X"08", X"f6", X"e5", X"0c", 
    X"24", X"f7", X"f8", X"e6", X"08", X"46", X"70", X"03", 
    X"02", X"55", X"c3", X"c0", X"e0", X"c0", X"a8", X"c2", 
    X"af", X"e5", X"0c", X"24", X"03", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"60", 
    X"56", X"aa", X"82", X"ab", X"83", X"e5", X"0c", X"24", 
    X"06", X"f8", X"a6", X"02", X"08", X"a6", X"03", X"e5", 
    X"0c", X"24", X"06", X"f8", X"e5", X"0c", X"24", X"08", 
    X"f9", X"c3", X"e7", X"96", X"09", X"e7", X"08", X"96", 
    X"92", X"00", X"40", X"4a", X"90", X"00", X"00", X"75", 
    X"f0", X"00", X"c0", X"20", X"12", X"21", X"e1", X"d0", 
    X"20", X"e5", X"0c", X"24", X"03", X"f8", X"74", X"08", 
    X"26", X"fa", X"e4", X"08", X"36", X"fb", X"08", X"86", 
    X"05", X"c0", X"05", X"c0", X"03", X"c0", X"02", X"c0", 
    X"20", X"12", X"15", X"47", X"ac", X"82", X"ae", X"83", 
    X"af", X"f0", X"d0", X"20", X"d0", X"02", X"d0", X"03", 
    X"d0", X"05", X"8a", X"82", X"8b", X"83", X"8d", X"f0", 
    X"ec", X"12", X"66", X"a0", X"a3", X"ee", X"12", X"66", 
    X"a0", X"a3", X"ef", X"12", X"66", X"a0", X"d0", X"e0", 
    X"53", X"e0", X"80", X"e5", X"e0", X"42", X"a8", X"d0", 
    X"e0", X"30", X"00", X"03", X"02", X"55", X"e1", X"e5", 
    X"0c", X"24", X"f7", X"f8", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"e4", X"c0", X"e0", X"c0", X"e0", 
    X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", 
    X"c0", X"e0", X"90", X"00", X"00", X"e4", X"f5", X"f0", 
    X"12", X"17", X"6d", X"e5", X"81", X"24", X"f7", X"f5", 
    X"81", X"e5", X"0c", X"24", X"03", X"f8", X"74", X"08", 
    X"26", X"fd", X"e4", X"08", X"36", X"fe", X"08", X"86", 
    X"07", X"7a", X"00", X"7b", X"00", X"7c", X"00", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"ea", X"12", X"66", 
    X"a0", X"a3", X"eb", X"12", X"66", X"a0", X"a3", X"ec", 
    X"12", X"66", X"a0", X"e5", X"0c", X"24", X"03", X"f8", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"12", X"60", X"56", X"ae", X"82", X"af", X"83", X"e5", 
    X"0c", X"24", X"06", X"f8", X"a6", X"06", X"08", X"a6", 
    X"07", X"80", X"1e", X"e5", X"0c", X"24", X"03", X"f8", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"12", X"60", X"56", X"ae", X"82", X"af", X"83", X"e5", 
    X"0c", X"24", X"06", X"f8", X"a6", X"06", X"08", X"a6", 
    X"07", X"e5", X"0c", X"24", X"06", X"f8", X"e5", X"0c", 
    X"24", X"08", X"f9", X"c3", X"e7", X"96", X"09", X"e7", 
    X"08", X"96", X"40", X"03", X"02", X"56", X"db", X"e5", 
    X"0c", X"24", X"08", X"f8", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"e5", X"0c", X"24", X"06", X"f8", 
    X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"e5", 
    X"0c", X"24", X"f9", X"f8", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"e5", X"0c", X"24", X"fb", X"f8", 
    X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"e5", X"0c", X"24", X"03", X"f8", 
    X"86", X"82", X"08", X"86", X"83", X"08", X"86", X"f0", 
    X"12", X"59", X"18", X"ae", X"82", X"af", X"83", X"e5", 
    X"81", X"24", X"f7", X"f5", X"81", X"a8", X"0c", X"08", 
    X"a6", X"06", X"08", X"a6", X"07", X"ee", X"4f", X"70", 
    X"03", X"02", X"56", X"db", X"12", X"09", X"4a", X"e5", 
    X"0c", X"24", X"03", X"f8", X"74", X"0b", X"26", X"fd", 
    X"e4", X"08", X"36", X"fe", X"08", X"86", X"07", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"fa", X"a3", X"12", X"70", X"5a", X"fb", X"a3", X"12", 
    X"70", X"5a", X"ea", X"4b", X"60", X"5a", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fa", 
    X"a3", X"12", X"70", X"5a", X"fb", X"a3", X"12", X"70", 
    X"5a", X"fc", X"c0", X"07", X"c0", X"06", X"c0", X"05", 
    X"e4", X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", 
    X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", 
    X"e0", X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"12", 
    X"19", X"e0", X"e5", X"81", X"24", X"f8", X"f5", X"81", 
    X"d0", X"05", X"d0", X"06", X"d0", X"07", X"7a", X"00", 
    X"7b", X"00", X"7c", X"00", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"ea", X"12", X"66", X"a0", X"a3", X"eb", 
    X"12", X"66", X"a0", X"a3", X"ec", X"12", X"66", X"a0", 
    X"12", X"09", X"52", X"a8", X"0c", X"08", X"86", X"82", 
    X"08", X"86", X"83", X"85", X"0c", X"81", X"d0", X"0c", 
    X"22", X"c0", X"0c", X"e5", X"81", X"f5", X"0c", X"24", 
    X"06", X"f5", X"81", X"ad", X"82", X"ae", X"83", X"af", 
    X"f0", X"74", X"11", X"2d", X"fa", X"e4", X"3e", X"fb", 
    X"8f", X"04", X"8a", X"82", X"8b", X"83", X"8c", X"f0", 
    X"12", X"70", X"5a", X"fa", X"20", X"e0", X"03", X"02", 
    X"57", X"b6", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"c0", X"07", X"c0", X"06", X"c0", X"05", X"12", X"60", 
    X"56", X"ab", X"82", X"ac", X"83", X"d0", X"05", X"d0", 
    X"06", X"d0", X"07", X"a8", X"0c", X"08", X"a6", X"03", 
    X"08", X"a6", X"04", X"a8", X"0c", X"08", X"c3", X"74", 
    X"02", X"96", X"e4", X"08", X"96", X"50", X"71", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"e5", X"0c", X"24", 
    X"03", X"f8", X"12", X"70", X"5a", X"f6", X"a3", X"12", 
    X"70", X"5a", X"08", X"f6", X"e5", X"0c", X"24", X"05", 
    X"fa", X"7b", X"00", X"7c", X"40", X"c0", X"07", X"c0", 
    X"06", X"c0", X"05", X"a8", X"0c", X"08", X"e6", X"c0", 
    X"e0", X"08", X"e6", X"c0", X"e0", X"74", X"02", X"c0", 
    X"e0", X"e4", X"c0", X"e0", X"c0", X"02", X"c0", X"03", 
    X"c0", X"04", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"12", X"5e", X"2e", X"e5", X"81", X"24", X"f9", X"f5", 
    X"81", X"d0", X"05", X"d0", X"06", X"d0", X"07", X"e5", 
    X"0c", X"24", X"05", X"f8", X"86", X"03", X"08", X"86", 
    X"04", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"e5", 
    X"0c", X"24", X"03", X"f8", X"e6", X"12", X"66", X"a0", 
    X"a3", X"08", X"e6", X"12", X"66", X"a0", X"80", X"0a", 
    X"7b", X"00", X"7c", X"00", X"80", X"04", X"7b", X"00", 
    X"7c", X"00", X"8b", X"82", X"8c", X"83", X"85", X"0c", 
    X"81", X"d0", X"0c", X"22", X"c0", X"0c", X"e5", X"81", 
    X"f5", X"0c", X"24", X"05", X"f5", X"81", X"af", X"82", 
    X"ae", X"83", X"ad", X"f0", X"e5", X"0c", X"24", X"03", 
    X"f8", X"a6", X"07", X"08", X"a6", X"06", X"08", X"a6", 
    X"05", X"a8", X"0c", X"08", X"e4", X"f6", X"08", X"f6", 
    X"74", X"11", X"2f", X"fb", X"e4", X"3e", X"fc", X"8b", 
    X"82", X"8c", X"83", X"8d", X"f0", X"12", X"70", X"5a", 
    X"30", X"e0", X"06", X"7c", X"02", X"7d", X"00", X"80", 
    X"04", X"7c", X"00", X"7d", X"00", X"e5", X"0c", X"24", 
    X"03", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"c0", X"05", X"c0", X"04", X"12", X"60", 
    X"56", X"aa", X"82", X"ab", X"83", X"d0", X"04", X"d0", 
    X"05", X"c3", X"ec", X"9a", X"ed", X"9b", X"40", X"03", 
    X"02", X"59", X"0a", X"c0", X"04", X"c0", X"05", X"c0", 
    X"02", X"c0", X"03", X"e5", X"0c", X"24", X"f9", X"f8", 
    X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"e5", 
    X"0c", X"24", X"fb", X"f8", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"e5", 
    X"0c", X"24", X"03", X"f8", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"59", X"18", X"ac", 
    X"82", X"ad", X"83", X"e5", X"81", X"24", X"f7", X"f5", 
    X"81", X"a8", X"0c", X"08", X"a6", X"04", X"08", X"a6", 
    X"05", X"ec", X"4d", X"70", X"03", X"02", X"59", X"0a", 
    X"e5", X"0c", X"24", X"03", X"f8", X"74", X"0b", X"26", 
    X"fb", X"e4", X"08", X"36", X"fc", X"08", X"86", X"05", 
    X"8b", X"82", X"8c", X"83", X"8d", X"f0", X"12", X"70", 
    X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"fe", X"a3", 
    X"12", X"70", X"5a", X"ff", X"ea", X"4e", X"60", X"6a", 
    X"8b", X"82", X"8c", X"83", X"8d", X"f0", X"12", X"70", 
    X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"fe", X"a3", 
    X"12", X"70", X"5a", X"ff", X"c0", X"05", X"c0", X"04", 
    X"c0", X"03", X"e5", X"0c", X"24", X"f6", X"f8", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"08", X"e6", 
    X"c0", X"e0", X"e4", X"c0", X"e0", X"c0", X"e0", X"c0", 
    X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", 
    X"e0", X"c0", X"e0", X"8a", X"82", X"8e", X"83", X"8f", 
    X"f0", X"12", X"1c", X"d7", X"e5", X"81", X"24", X"f5", 
    X"f5", X"81", X"d0", X"03", X"d0", X"04", X"d0", X"05", 
    X"7a", X"00", X"7e", X"00", X"7f", X"00", X"8b", X"82", 
    X"8c", X"83", X"8d", X"f0", X"ea", X"12", X"66", X"a0", 
    X"a3", X"ee", X"12", X"66", X"a0", X"a3", X"ef", X"12", 
    X"66", X"a0", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"85", X"0c", X"81", X"d0", X"0c", X"22", 
    X"c0", X"0c", X"e5", X"81", X"f5", X"0c", X"24", X"06", 
    X"f5", X"81", X"ad", X"82", X"ae", X"83", X"af", X"f0", 
    X"e5", X"0c", X"24", X"f5", X"f8", X"e6", X"08", X"46", 
    X"70", X"03", X"02", X"59", X"de", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"a8", X"0c", X"08", X"12", X"70", 
    X"5a", X"f6", X"a3", X"12", X"70", X"5a", X"08", X"f6", 
    X"e5", X"0c", X"24", X"05", X"fa", X"7b", X"00", X"7c", 
    X"40", X"c0", X"07", X"c0", X"06", X"c0", X"05", X"e5", 
    X"0c", X"24", X"f7", X"f8", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"e5", X"0c", X"24", X"f5", X"f8", 
    X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"c0", 
    X"02", X"c0", X"03", X"c0", X"04", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"5e", X"2e", X"e5", X"81", 
    X"24", X"f9", X"f5", X"81", X"d0", X"05", X"d0", X"06", 
    X"d0", X"07", X"e5", X"0c", X"24", X"05", X"f8", X"e5", 
    X"0c", X"24", X"03", X"f9", X"e6", X"f7", X"08", X"09", 
    X"e6", X"f7", X"e5", X"0c", X"24", X"f7", X"f8", X"e5", 
    X"0c", X"24", X"f5", X"f9", X"e6", X"c3", X"97", X"f6", 
    X"08", X"e6", X"09", X"97", X"f6", X"e5", X"0c", X"24", 
    X"03", X"f8", X"e5", X"0c", X"24", X"f9", X"f9", X"c3", 
    X"e7", X"96", X"09", X"e7", X"08", X"96", X"50", X"2e", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"a8", X"0c", 
    X"08", X"e6", X"12", X"66", X"a0", X"a3", X"08", X"e6", 
    X"12", X"66", X"a0", X"e5", X"0c", X"24", X"03", X"f8", 
    X"e4", X"f6", X"08", X"f6", X"80", X"10", X"e5", X"0c", 
    X"24", X"f9", X"f8", X"e5", X"0c", X"24", X"03", X"f9", 
    X"e6", X"f7", X"08", X"09", X"e6", X"f7", X"e5", X"0c", 
    X"24", X"fb", X"f8", X"86", X"02", X"08", X"86", X"03", 
    X"08", X"86", X"04", X"e5", X"0c", X"24", X"f7", X"f8", 
    X"e6", X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"e5", 
    X"0c", X"24", X"03", X"f8", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"c0", X"02", X"c0", X"03", X"c0", 
    X"04", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"5e", X"2e", X"ae", X"82", X"af", X"83", X"e5", X"81", 
    X"24", X"f9", X"f5", X"81", X"8e", X"82", X"8f", X"83", 
    X"85", X"0c", X"81", X"d0", X"0c", X"22", X"ad", X"82", 
    X"ae", X"83", X"af", X"f0", X"12", X"70", X"5a", X"fb", 
    X"a3", X"12", X"70", X"5a", X"fc", X"74", X"02", X"2d", 
    X"fd", X"e4", X"3e", X"fe", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"70", X"5a", X"fd", X"a3", X"12", 
    X"70", X"5a", X"fe", X"ed", X"b5", X"03", X"08", X"ee", 
    X"b5", X"04", X"04", X"7f", X"01", X"80", X"02", X"7f", 
    X"00", X"8f", X"82", X"22", X"ad", X"82", X"ae", X"83", 
    X"af", X"f0", X"74", X"11", X"2d", X"fa", X"e4", X"3e", 
    X"fb", X"8f", X"04", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"12", X"70", X"5a", X"30", X"e0", X"06", X"7b", 
    X"02", X"7c", X"00", X"80", X"04", X"7b", X"00", X"7c", 
    X"00", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"c0", 
    X"04", X"c0", X"03", X"12", X"4e", X"60", X"ae", X"82", 
    X"af", X"83", X"d0", X"03", X"d0", X"04", X"c3", X"eb", 
    X"9e", X"ec", X"9f", X"40", X"04", X"7f", X"01", X"80", 
    X"02", X"7f", X"00", X"8f", X"82", X"22", X"c0", X"0c", 
    X"85", X"81", X"0c", X"ad", X"82", X"ae", X"83", X"af", 
    X"f0", X"74", X"08", X"2d", X"fd", X"e4", X"3e", X"fe", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", 
    X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"fb", X"a3", 
    X"12", X"70", X"5a", X"fc", X"ea", X"4b", X"60", X"6e", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", 
    X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"fb", X"a3", 
    X"12", X"70", X"5a", X"fc", X"c0", X"07", X"c0", X"06", 
    X"c0", X"05", X"e5", X"0c", X"24", X"fb", X"f8", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"08", X"e6", 
    X"c0", X"e0", X"e4", X"c0", X"e0", X"c0", X"e0", X"c0", 
    X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", 
    X"e0", X"c0", X"e0", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"12", X"1c", X"d7", X"e5", X"81", X"24", X"f5", 
    X"f5", X"81", X"d0", X"05", X"d0", X"06", X"d0", X"07", 
    X"7a", X"00", X"7b", X"00", X"7c", X"00", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"ea", X"12", X"66", X"a0", 
    X"a3", X"eb", X"12", X"66", X"a0", X"a3", X"ec", X"12", 
    X"66", X"a0", X"7f", X"01", X"80", X"02", X"7f", X"00", 
    X"8f", X"82", X"d0", X"0c", X"22", X"c0", X"0c", X"85", 
    X"81", X"0c", X"ad", X"82", X"ae", X"83", X"af", X"f0", 
    X"74", X"0b", X"2d", X"fd", X"e4", X"3e", X"fe", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"fa", X"a3", X"12", X"70", X"5a", X"fb", X"a3", X"12", 
    X"70", X"5a", X"fc", X"ea", X"4b", X"60", X"6e", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"fa", X"a3", X"12", X"70", X"5a", X"fb", X"a3", X"12", 
    X"70", X"5a", X"fc", X"c0", X"07", X"c0", X"06", X"c0", 
    X"05", X"e5", X"0c", X"24", X"fb", X"f8", X"e6", X"c0", 
    X"e0", X"08", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"e4", X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", 
    X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", X"c0", X"e0", 
    X"c0", X"e0", X"8a", X"82", X"8b", X"83", X"8c", X"f0", 
    X"12", X"1c", X"d7", X"e5", X"81", X"24", X"f5", X"f5", 
    X"81", X"d0", X"05", X"d0", X"06", X"d0", X"07", X"7a", 
    X"00", X"7b", X"00", X"7c", X"00", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"ea", X"12", X"66", X"a0", X"a3", 
    X"eb", X"12", X"66", X"a0", X"a3", X"ec", X"12", X"66", 
    X"a0", X"7f", X"01", X"80", X"02", X"7f", X"00", X"8f", 
    X"82", X"d0", X"0c", X"22", X"c0", X"0c", X"85", X"81", 
    X"0c", X"c0", X"82", X"c0", X"83", X"c0", X"f0", X"e5", 
    X"81", X"24", X"0c", X"f5", X"81", X"a8", X"0c", X"08", 
    X"74", X"02", X"26", X"fa", X"e4", X"08", X"36", X"fb", 
    X"08", X"86", X"04", X"8a", X"82", X"8b", X"83", X"8c", 
    X"f0", X"e5", X"0c", X"24", X"04", X"f8", X"12", X"70", 
    X"5a", X"f6", X"a3", X"12", X"70", X"5a", X"08", X"f6", 
    X"a8", X"0c", X"08", X"e5", X"0c", X"24", X"06", X"f9", 
    X"74", X"04", X"26", X"f7", X"e4", X"08", X"36", X"09", 
    X"f7", X"08", X"09", X"e6", X"f7", X"e5", X"0c", X"24", 
    X"06", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"e5", X"0c", X"24", X"09", X"f9", X"12", 
    X"70", X"5a", X"f7", X"a3", X"12", X"70", X"5a", X"09", 
    X"f7", X"e5", X"0c", X"24", X"09", X"f8", X"e5", X"0c", 
    X"24", X"04", X"f9", X"e6", X"c3", X"97", X"fe", X"08", 
    X"e6", X"09", X"97", X"ff", X"e5", X"0c", X"24", X"f9", 
    X"f8", X"c3", X"ee", X"96", X"ef", X"08", X"96", X"50", 
    X"15", X"e5", X"0c", X"24", X"09", X"f8", X"e5", X"0c", 
    X"24", X"04", X"f9", X"e6", X"c3", X"97", X"fe", X"08", 
    X"e6", X"09", X"97", X"ff", X"80", X"0a", X"e5", X"0c", 
    X"24", X"f9", X"f8", X"86", X"06", X"08", X"86", X"07", 
    X"c0", X"02", X"c0", X"03", X"c0", X"04", X"e5", X"0c", 
    X"24", X"0e", X"f8", X"a6", X"06", X"08", X"a6", X"07", 
    X"e5", X"0c", X"24", X"fb", X"f8", X"86", X"03", X"08", 
    X"86", X"04", X"08", X"86", X"05", X"a8", X"0c", X"08", 
    X"e5", X"0c", X"24", X"0b", X"f9", X"74", X"0e", X"26", 
    X"f7", X"e4", X"08", X"36", X"09", X"f7", X"08", X"09", 
    X"e6", X"f7", X"e5", X"0c", X"24", X"0b", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"12", 
    X"70", X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"fe", 
    X"a3", X"12", X"70", X"5a", X"ff", X"e5", X"0c", X"24", 
    X"04", X"f8", X"e6", X"2a", X"fa", X"08", X"e6", X"3e", 
    X"fe", X"c0", X"04", X"c0", X"03", X"c0", X"02", X"e5", 
    X"0c", X"24", X"0e", X"f8", X"e6", X"c0", X"e0", X"08", 
    X"e6", X"c0", X"e0", X"c0", X"03", X"c0", X"04", X"c0", 
    X"05", X"8a", X"82", X"8e", X"83", X"8f", X"f0", X"12", 
    X"67", X"03", X"e5", X"81", X"24", X"fb", X"f5", X"81", 
    X"d0", X"02", X"d0", X"03", X"d0", X"04", X"e5", X"0c", 
    X"24", X"f9", X"f8", X"e5", X"0c", X"24", X"0e", X"f9", 
    X"c3", X"e7", X"96", X"09", X"e7", X"08", X"96", X"d0", 
    X"04", X"d0", X"03", X"d0", X"02", X"40", X"03", X"02", 
    X"5d", X"c7", X"c0", X"02", X"c0", X"03", X"c0", X"04", 
    X"e5", X"0c", X"24", X"f9", X"f8", X"e5", X"0c", X"24", 
    X"0e", X"f9", X"e6", X"c3", X"97", X"c0", X"e0", X"08", 
    X"e6", X"09", X"97", X"c0", X"e0", X"e5", X"0c", X"24", 
    X"0a", X"f8", X"d0", X"e0", X"f6", X"18", X"d0", X"e0", 
    X"f6", X"e5", X"0c", X"24", X"fb", X"f8", X"e5", X"0c", 
    X"24", X"0e", X"f9", X"e7", X"26", X"fb", X"09", X"e7", 
    X"08", X"36", X"08", X"86", X"05", X"7d", X"00", X"7c", 
    X"40", X"e5", X"0c", X"24", X"0b", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"12", X"70", 
    X"5a", X"fa", X"a3", X"12", X"70", X"5a", X"fe", X"a3", 
    X"12", X"70", X"5a", X"ff", X"c0", X"04", X"c0", X"03", 
    X"c0", X"02", X"e5", X"0c", X"24", X"09", X"f8", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"c0", X"03", 
    X"c0", X"05", X"c0", X"04", X"8a", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"67", X"03", X"e5", X"81", X"24", 
    X"fb", X"f5", X"81", X"d0", X"02", X"d0", X"03", X"d0", 
    X"04", X"d0", X"04", X"d0", X"03", X"d0", X"02", X"e5", 
    X"0c", X"24", X"04", X"f8", X"e5", X"0c", X"24", X"f9", 
    X"f9", X"e7", X"26", X"fe", X"09", X"e7", X"08", X"36", 
    X"ff", X"e5", X"0c", X"24", X"06", X"f8", X"86", X"82", 
    X"08", X"86", X"83", X"08", X"86", X"f0", X"e5", X"0c", 
    X"24", X"0b", X"f9", X"12", X"70", X"5a", X"f7", X"a3", 
    X"12", X"70", X"5a", X"09", X"f7", X"e5", X"0c", X"24", 
    X"0b", X"f8", X"c3", X"ee", X"96", X"ef", X"08", X"96", 
    X"40", X"0d", X"e5", X"0c", X"24", X"0b", X"f8", X"ee", 
    X"c3", X"96", X"fe", X"ef", X"08", X"96", X"ff", X"8a", 
    X"82", X"8b", X"83", X"8c", X"f0", X"ee", X"12", X"66", 
    X"a0", X"a3", X"ef", X"12", X"66", X"a0", X"e5", X"0c", 
    X"24", X"f9", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"85", X"0c", X"81", X"d0", X"0c", X"22", X"c0", X"0c", 
    X"85", X"81", X"0c", X"c0", X"82", X"c0", X"83", X"c0", 
    X"f0", X"e5", X"81", X"24", X"0c", X"f5", X"81", X"e5", 
    X"0c", X"24", X"f7", X"f8", X"e5", X"0c", X"24", X"f9", 
    X"f9", X"c3", X"e6", X"97", X"08", X"e6", X"09", X"97", 
    X"50", X"0c", X"e5", X"0c", X"24", X"f7", X"f8", X"86", 
    X"03", X"08", X"86", X"04", X"80", X"0a", X"e5", X"0c", 
    X"24", X"f9", X"f8", X"86", X"03", X"08", X"86", X"04", 
    X"e5", X"0c", X"24", X"0c", X"f8", X"a6", X"03", X"08", 
    X"a6", X"04", X"e5", X"0c", X"24", X"0c", X"f8", X"e6", 
    X"08", X"46", X"70", X"03", X"02", X"60", X"46", X"a8", 
    X"0c", X"08", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"12", X"70", X"5a", X"fa", X"a3", X"12", 
    X"70", X"5a", X"fc", X"a8", X"0c", X"08", X"e5", X"0c", 
    X"24", X"04", X"f9", X"74", X"04", X"26", X"f7", X"e4", 
    X"08", X"36", X"09", X"f7", X"08", X"09", X"e6", X"f7", 
    X"e5", X"0c", X"24", X"04", X"f8", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", 
    X"fe", X"a3", X"12", X"70", X"5a", X"fd", X"ee", X"c3", 
    X"9a", X"fb", X"ed", X"9c", X"ff", X"e5", X"0c", X"24", 
    X"0c", X"f8", X"c3", X"eb", X"96", X"ef", X"08", X"96", 
    X"50", X"09", X"ee", X"c3", X"9a", X"fe", X"ed", X"9c", 
    X"ff", X"80", X"0a", X"e5", X"0c", X"24", X"0c", X"f8", 
    X"86", X"06", X"08", X"86", X"07", X"e5", X"0c", X"24", 
    X"0e", X"f8", X"a6", X"06", X"08", X"a6", X"07", X"a8", 
    X"0c", X"08", X"e5", X"0c", X"24", X"09", X"f9", X"74", 
    X"0e", X"26", X"f7", X"e4", X"08", X"36", X"09", X"f7", 
    X"08", X"09", X"e6", X"f7", X"e5", X"0c", X"24", X"09", 
    X"f8", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"12", X"70", X"5a", X"fd", X"a3", X"12", X"70", 
    X"5a", X"fe", X"a3", X"12", X"70", X"5a", X"ff", X"ea", 
    X"2d", X"fd", X"ec", X"3e", X"fe", X"c0", X"02", X"c0", 
    X"04", X"e5", X"0c", X"24", X"fb", X"f8", X"86", X"02", 
    X"08", X"86", X"03", X"08", X"86", X"04", X"c0", X"04", 
    X"c0", X"02", X"e5", X"0c", X"24", X"0e", X"f8", X"e6", 
    X"c0", X"e0", X"08", X"e6", X"c0", X"e0", X"c0", X"05", 
    X"c0", X"06", X"c0", X"07", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"12", X"67", X"03", X"e5", X"81", X"24", 
    X"fb", X"f5", X"81", X"d0", X"02", X"d0", X"04", X"e5", 
    X"0c", X"24", X"0c", X"f8", X"e5", X"0c", X"24", X"0e", 
    X"f9", X"c3", X"e7", X"96", X"09", X"e7", X"08", X"96", 
    X"d0", X"04", X"d0", X"02", X"40", X"03", X"02", X"5f", 
    X"fe", X"c0", X"02", X"c0", X"04", X"e5", X"0c", X"24", 
    X"0c", X"f8", X"e5", X"0c", X"24", X"0e", X"f9", X"e6", 
    X"c3", X"97", X"c0", X"e0", X"08", X"e6", X"09", X"97", 
    X"c0", X"e0", X"e5", X"0c", X"24", X"08", X"f8", X"d0", 
    X"e0", X"f6", X"18", X"d0", X"e0", X"f6", X"e5", X"0c", 
    X"24", X"09", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"70", X"5a", X"fb", X"a3", 
    X"12", X"70", X"5a", X"fc", X"a3", X"12", X"70", X"5a", 
    X"fd", X"e5", X"0c", X"24", X"fb", X"f8", X"e5", X"0c", 
    X"24", X"0e", X"f9", X"e7", X"26", X"fa", X"09", X"e7", 
    X"08", X"36", X"08", X"86", X"07", X"7f", X"00", X"7e", 
    X"40", X"c0", X"04", X"c0", X"02", X"e5", X"0c", X"24", 
    X"07", X"f8", X"e6", X"c0", X"e0", X"08", X"e6", X"c0", 
    X"e0", X"c0", X"03", X"c0", X"04", X"c0", X"05", X"8a", 
    X"82", X"8f", X"83", X"8e", X"f0", X"12", X"67", X"03", 
    X"e5", X"81", X"24", X"fb", X"f5", X"81", X"d0", X"02", 
    X"d0", X"04", X"d0", X"04", X"d0", X"02", X"e5", X"0c", 
    X"24", X"0c", X"f8", X"e6", X"2a", X"fa", X"08", X"e6", 
    X"3c", X"fc", X"8a", X"07", X"8c", X"06", X"e5", X"0c", 
    X"24", X"04", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"12", X"70", X"5a", X"fc", X"a3", 
    X"12", X"70", X"5a", X"fd", X"c3", X"ef", X"9c", X"ee", 
    X"9d", X"40", X"07", X"ef", X"c3", X"9c", X"ff", X"ee", 
    X"9d", X"fe", X"a8", X"0c", X"08", X"86", X"82", X"08", 
    X"86", X"83", X"08", X"86", X"f0", X"ef", X"12", X"66", 
    X"a0", X"a3", X"ee", X"12", X"66", X"a0", X"e5", X"0c", 
    X"24", X"0c", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"85", X"0c", X"81", X"d0", X"0c", X"22", X"c0", X"0c", 
    X"85", X"81", X"0c", X"c0", X"82", X"c0", X"83", X"c0", 
    X"f0", X"a8", X"0c", X"08", X"74", X"04", X"26", X"fb", 
    X"e4", X"08", X"36", X"fa", X"08", X"86", X"04", X"8b", 
    X"82", X"8a", X"83", X"8c", X"f0", X"12", X"70", X"5a", 
    X"fb", X"a3", X"12", X"70", X"5a", X"fc", X"a8", X"0c", 
    X"08", X"74", X"02", X"26", X"fa", X"e4", X"08", X"36", 
    X"fe", X"08", X"86", X"07", X"8a", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"70", X"5a", X"fa", X"a3", X"12", 
    X"70", X"5a", X"fe", X"ea", X"2b", X"fa", X"ee", X"3c", 
    X"fe", X"a8", X"0c", X"08", X"86", X"82", X"08", X"86", 
    X"83", X"08", X"86", X"f0", X"12", X"70", X"5a", X"fd", 
    X"a3", X"12", X"70", X"5a", X"ff", X"ea", X"c3", X"9d", 
    X"fd", X"ee", X"9f", X"ff", X"8d", X"06", X"c3", X"ee", 
    X"9b", X"ef", X"9c", X"40", X"07", X"ee", X"c3", X"9b", 
    X"fe", X"ef", X"9c", X"ff", X"8e", X"82", X"8f", X"83", 
    X"85", X"0c", X"81", X"d0", X"0c", X"22", X"c0", X"0c", 
    X"85", X"81", X"0c", X"ad", X"82", X"ae", X"83", X"af", 
    X"f0", X"8d", X"02", X"8e", X"03", X"8f", X"04", X"c0", 
    X"07", X"c0", X"06", X"c0", X"05", X"74", X"12", X"c0", 
    X"e0", X"e4", X"c0", X"e0", X"c0", X"e0", X"8a", X"82", 
    X"8b", X"83", X"8c", X"f0", X"12", X"66", X"db", X"15", 
    X"81", X"15", X"81", X"15", X"81", X"d0", X"05", X"d0", 
    X"06", X"d0", X"07", X"74", X"0e", X"2d", X"fa", X"e4", 
    X"3e", X"fb", X"8f", X"04", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"e5", X"0c", X"24", X"fb", X"f8", X"e6", 
    X"12", X"66", X"a0", X"a3", X"08", X"e6", X"12", X"66", 
    X"a0", X"a3", X"08", X"e6", X"12", X"66", X"a0", X"74", 
    X"04", X"2d", X"fa", X"e4", X"3e", X"fb", X"8f", X"04", 
    X"8a", X"82", X"8b", X"83", X"8c", X"f0", X"e5", X"0c", 
    X"24", X"f9", X"f8", X"e6", X"12", X"66", X"a0", X"a3", 
    X"08", X"e6", X"12", X"66", X"a0", X"74", X"06", X"2d", 
    X"fa", X"e4", X"3e", X"fb", X"8f", X"04", X"8a", X"82", 
    X"8b", X"83", X"8c", X"f0", X"e5", X"0c", X"24", X"f7", 
    X"f8", X"e6", X"12", X"66", X"a0", X"a3", X"08", X"e6", 
    X"12", X"66", X"a0", X"74", X"11", X"2d", X"fd", X"e4", 
    X"3e", X"fe", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"e5", X"0c", X"24", X"f6", X"f8", X"e6", X"12", X"66", 
    X"a0", X"d0", X"0c", X"22", X"c0", X"0c", X"85", X"81", 
    X"0c", X"c0", X"82", X"c0", X"83", X"05", X"81", X"05", 
    X"81", X"05", X"81", X"e5", X"0c", X"24", X"03", X"f8", 
    X"e4", X"f6", X"08", X"f6", X"08", X"76", X"00", X"12", 
    X"09", X"4a", X"90", X"18", X"77", X"e0", X"f5", X"f0", 
    X"a3", X"e0", X"45", X"f0", X"70", X"11", X"7a", X"76", 
    X"7d", X"00", X"fe", X"ff", X"90", X"18", X"77", X"ea", 
    X"f0", X"ed", X"a3", X"f0", X"ee", X"a3", X"f0", X"90", 
    X"18", X"75", X"e0", X"fe", X"a3", X"e0", X"ff", X"a8", 
    X"0c", X"08", X"e6", X"2e", X"fc", X"08", X"e6", X"3f", 
    X"fd", X"c3", X"ec", X"94", X"ff", X"ed", X"94", X"17", 
    X"50", X"3d", X"a8", X"0c", X"08", X"e6", X"2e", X"fc", 
    X"08", X"e6", X"3f", X"fd", X"c3", X"ee", X"9c", X"ef", 
    X"9d", X"50", X"2c", X"90", X"18", X"77", X"e0", X"fb", 
    X"a3", X"e0", X"fc", X"a3", X"e0", X"fd", X"ee", X"2b", 
    X"fb", X"ef", X"3c", X"fc", X"e5", X"0c", X"24", X"03", 
    X"f8", X"a6", X"03", X"08", X"a6", X"04", X"08", X"a6", 
    X"05", X"a8", X"0c", X"08", X"90", X"18", X"75", X"e6", 
    X"2e", X"f0", X"08", X"e6", X"3f", X"a3", X"f0", X"12", 
    X"09", X"52", X"e5", X"0c", X"24", X"03", X"f8", X"86", 
    X"82", X"08", X"86", X"83", X"08", X"86", X"f0", X"85", 
    X"0c", X"81", X"d0", X"0c", X"22", X"22", X"90", X"18", 
    X"75", X"e4", X"f0", X"a3", X"f0", X"22", X"90", X"18", 
    X"75", X"e0", X"fe", X"a3", X"e0", X"ff", X"74", X"ff", 
    X"c3", X"9e", X"fe", X"74", X"17", X"9f", X"8e", X"82", 
    X"f5", X"83", X"22", X"c0", X"0c", X"e5", X"81", X"f5", 
    X"0c", X"24", X"0e", X"f5", X"81", X"ad", X"82", X"ae", 
    X"83", X"af", X"f0", X"e5", X"0c", X"24", X"0c", X"f8", 
    X"a6", X"05", X"08", X"a6", X"06", X"08", X"a6", X"07", 
    X"a8", X"0c", X"08", X"74", X"01", X"2d", X"f6", X"e4", 
    X"3e", X"08", X"f6", X"08", X"a6", X"07", X"e5", X"0c", 
    X"24", X"fc", X"f8", X"86", X"02", X"08", X"86", X"03", 
    X"7c", X"80", X"7f", X"00", X"8a", X"06", X"a8", X"0c", 
    X"08", X"86", X"82", X"08", X"86", X"83", X"08", X"86", 
    X"f0", X"ee", X"12", X"66", X"a0", X"e5", X"0c", X"24", 
    X"04", X"f8", X"a6", X"03", X"08", X"a6", X"04", X"08", 
    X"a6", X"07", X"08", X"76", X"00", X"a8", X"0c", X"08", 
    X"74", X"01", X"26", X"fd", X"e4", X"08", X"36", X"fe", 
    X"08", X"86", X"07", X"e5", X"0c", X"24", X"04", X"f8", 
    X"86", X"02", X"8d", X"82", X"8e", X"83", X"8f", X"f0", 
    X"ea", X"12", X"66", X"a0", X"0d", X"bd", X"00", X"01", 
    X"0e", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"74", 
    X"aa", X"12", X"66", X"a0", X"0d", X"bd", X"00", X"01", 
    X"0e", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"74", 
    X"80", X"12", X"66", X"a0", X"e5", X"0c", X"24", X"04", 
    X"f8", X"74", X"01", X"2d", X"f6", X"e4", X"3e", X"08", 
    X"f6", X"08", X"a6", X"07", X"e5", X"0c", X"24", X"f9", 
    X"f8", X"86", X"02", X"08", X"86", X"03", X"08", X"86", 
    X"04", X"7f", X"00", X"8a", X"06", X"e5", X"0c", X"24", 
    X"04", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"ee", X"12", X"66", X"a0", X"e5", X"0c", 
    X"24", X"08", X"f8", X"a6", X"03", X"08", X"a6", X"04", 
    X"08", X"a6", X"07", X"08", X"76", X"00", X"e5", X"0c", 
    X"24", X"04", X"f8", X"74", X"01", X"26", X"fd", X"e4", 
    X"08", X"36", X"fe", X"08", X"86", X"07", X"e5", X"0c", 
    X"24", X"08", X"f8", X"86", X"02", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"ea", X"12", X"66", X"a0", X"e5", 
    X"0c", X"24", X"08", X"f8", X"08", X"e6", X"18", X"f6", 
    X"08", X"08", X"e6", X"18", X"f6", X"08", X"08", X"e6", 
    X"18", X"f6", X"08", X"76", X"00", X"0d", X"bd", X"00", 
    X"01", X"0e", X"e5", X"0c", X"24", X"08", X"f8", X"86", 
    X"02", X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"ea", 
    X"12", X"66", X"a0", X"0d", X"bd", X"00", X"01", X"0e", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"74", X"02", 
    X"12", X"66", X"a0", X"0d", X"bd", X"00", X"01", X"0e", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"74", X"03", 
    X"12", X"66", X"a0", X"0d", X"bd", X"00", X"01", X"0e", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"74", X"04", 
    X"12", X"66", X"a0", X"0d", X"bd", X"00", X"01", X"0e", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"74", X"05", 
    X"12", X"66", X"a0", X"0d", X"bd", X"00", X"01", X"0e", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"74", X"06", 
    X"12", X"66", X"a0", X"0d", X"bd", X"00", X"01", X"0e", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"74", X"07", 
    X"12", X"66", X"a0", X"0d", X"bd", X"00", X"01", X"0e", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"e4", X"12", 
    X"66", X"a0", X"0d", X"bd", X"00", X"01", X"0e", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"74", X"01", X"12", 
    X"66", X"a0", X"0d", X"bd", X"00", X"01", X"0e", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"e4", X"12", X"66", 
    X"a0", X"0d", X"bd", X"00", X"01", X"0e", X"8d", X"82", 
    X"8e", X"83", X"8f", X"f0", X"74", X"bb", X"12", X"66", 
    X"a0", X"e5", X"0c", X"24", X"0c", X"f8", X"ed", X"c3", 
    X"96", X"fd", X"ee", X"08", X"96", X"e5", X"0c", X"24", 
    X"0c", X"f8", X"86", X"82", X"08", X"86", X"83", X"08", 
    X"86", X"f0", X"ed", X"12", X"66", X"a0", X"e5", X"0c", 
    X"24", X"0c", X"f8", X"86", X"82", X"08", X"86", X"83", 
    X"08", X"86", X"f0", X"85", X"0c", X"81", X"d0", X"0c", 
    X"22", X"12", X"66", X"76", X"90", X"00", X"09", X"e0", 
    X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"f5", X"09", X"a3", X"12", X"70", X"5a", X"f5", X"0a", 
    X"75", X"0b", X"0d", X"85", X"09", X"82", X"85", X"0a", 
    X"83", X"e0", X"f5", X"08", X"05", X"09", X"e4", X"b5", 
    X"09", X"02", X"05", X"0a", X"05", X"0b", X"a9", X"0b", 
    X"85", X"09", X"82", X"85", X"0a", X"83", X"e0", X"ff", 
    X"f7", X"d5", X"08", X"e8", X"85", X"0b", X"81", X"d0", 
    X"0c", X"d0", X"d0", X"d0", X"01", X"d0", X"00", X"d0", 
    X"07", X"d0", X"06", X"d0", X"05", X"d0", X"04", X"d0", 
    X"03", X"d0", X"02", X"d0", X"f0", X"d0", X"83", X"d0", 
    X"82", X"d0", X"e0", X"20", X"e7", X"05", X"c2", X"af", 
    X"02", X"64", X"ad", X"d2", X"af", X"d0", X"e0", X"32", 
    X"75", X"82", X"01", X"22", X"22", X"c0", X"e0", X"c0", 
    X"a8", X"c2", X"af", X"c0", X"82", X"c0", X"83", X"c0", 
    X"f0", X"c0", X"02", X"c0", X"03", X"c0", X"04", X"c0", 
    X"05", X"c0", X"06", X"c0", X"07", X"c0", X"00", X"c0", 
    X"01", X"c0", X"d0", X"75", X"d0", X"00", X"c0", X"0c", 
    X"90", X"00", X"09", X"e0", X"fd", X"a3", X"e0", X"fe", 
    X"a3", X"e0", X"ff", X"8d", X"82", X"8e", X"83", X"8f", 
    X"f0", X"12", X"70", X"5a", X"f5", X"09", X"a3", X"12", 
    X"70", X"5a", X"f5", X"0a", X"75", X"0b", X"0e", X"e5", 
    X"81", X"ff", X"24", X"f3", X"f5", X"08", X"85", X"09", 
    X"82", X"85", X"0a", X"83", X"f0", X"e5", X"08", X"60", 
    X"19", X"05", X"09", X"e4", X"b5", X"09", X"02", X"05", 
    X"0a", X"85", X"09", X"82", X"85", X"0a", X"83", X"a9", 
    X"0b", X"e7", X"ff", X"f0", X"05", X"0b", X"15", X"08", 
    X"80", X"e3", X"12", X"0e", X"13", X"90", X"00", X"09", 
    X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", 
    X"5a", X"f5", X"09", X"a3", X"12", X"70", X"5a", X"f5", 
    X"0a", X"75", X"0b", X"0d", X"85", X"09", X"82", X"85", 
    X"0a", X"83", X"e0", X"f5", X"08", X"05", X"09", X"e4", 
    X"b5", X"09", X"02", X"05", X"0a", X"05", X"0b", X"a9", 
    X"0b", X"85", X"09", X"82", X"85", X"0a", X"83", X"e0", 
    X"ff", X"f7", X"d5", X"08", X"e8", X"85", X"0b", X"81", 
    X"d0", X"0c", X"d0", X"d0", X"d0", X"01", X"d0", X"00", 
    X"d0", X"07", X"d0", X"06", X"d0", X"05", X"d0", X"04", 
    X"d0", X"03", X"d0", X"02", X"d0", X"f0", X"d0", X"83", 
    X"d0", X"82", X"d0", X"e0", X"20", X"e7", X"05", X"c2", 
    X"af", X"02", X"65", X"8e", X"d2", X"af", X"d0", X"e0", 
    X"32", X"c0", X"e0", X"c0", X"a8", X"c2", X"af", X"c0", 
    X"82", X"c0", X"83", X"c0", X"f0", X"c0", X"02", X"c0", 
    X"03", X"c0", X"04", X"c0", X"05", X"c0", X"06", X"c0", 
    X"07", X"c0", X"00", X"c0", X"01", X"c0", X"d0", X"75", 
    X"d0", X"00", X"c0", X"0c", X"90", X"00", X"09", X"e0", 
    X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"f5", X"09", X"a3", X"12", X"70", X"5a", X"f5", X"0a", 
    X"75", X"0b", X"0e", X"e5", X"81", X"ff", X"24", X"f3", 
    X"f5", X"08", X"85", X"09", X"82", X"85", X"0a", X"83", 
    X"f0", X"e5", X"08", X"60", X"19", X"05", X"09", X"e4", 
    X"b5", X"09", X"02", X"05", X"0a", X"85", X"09", X"82", 
    X"85", X"0a", X"83", X"a9", X"0b", X"e7", X"ff", X"f0", 
    X"05", X"0b", X"15", X"08", X"80", X"e3", X"12", X"0b", 
    X"66", X"e5", X"82", X"60", X"03", X"12", X"0e", X"13", 
    X"d2", X"88", X"90", X"00", X"09", X"e0", X"fd", X"a3", 
    X"e0", X"fe", X"a3", X"e0", X"ff", X"8d", X"82", X"8e", 
    X"83", X"8f", X"f0", X"12", X"70", X"5a", X"f5", X"09", 
    X"a3", X"12", X"70", X"5a", X"f5", X"0a", X"75", X"0b", 
    X"0d", X"85", X"09", X"82", X"85", X"0a", X"83", X"e0", 
    X"f5", X"08", X"05", X"09", X"e4", X"b5", X"09", X"02", 
    X"05", X"0a", X"05", X"0b", X"a9", X"0b", X"85", X"09", 
    X"82", X"85", X"0a", X"83", X"e0", X"ff", X"f7", X"d5", 
    X"08", X"e8", X"85", X"0b", X"81", X"d0", X"0c", X"d0", 
    X"d0", X"d0", X"01", X"d0", X"00", X"d0", X"07", X"d0", 
    X"06", X"d0", X"05", X"d0", X"04", X"d0", X"03", X"d0", 
    X"02", X"d0", X"f0", X"d0", X"83", X"d0", X"82", X"d0", 
    X"e0", X"20", X"e7", X"05", X"c2", X"af", X"02", X"66", 
    X"73", X"d2", X"af", X"d0", X"e0", X"32", X"75", X"8f", 
    X"fc", X"75", X"8e", X"18", X"d2", X"8c", X"d2", X"88", 
    X"d2", X"a9", X"d2", X"af", X"d2", X"8d", X"22", X"af", 
    X"82", X"30", X"9c", X"fd", X"8f", X"99", X"bf", X"0a", 
    X"06", X"30", X"9c", X"fd", X"75", X"99", X"0d", X"22", 
    X"30", X"9d", X"fd", X"af", X"99", X"8f", X"82", X"22", 
    X"20", X"f7", X"11", X"30", X"f6", X"13", X"88", X"83", 
    X"a8", X"82", X"20", X"f5", X"09", X"f6", X"a8", X"83", 
    X"75", X"83", X"00", X"22", X"80", X"fe", X"f2", X"80", 
    X"f5", X"f0", X"22", X"aa", X"83", X"ab", X"82", X"8b", 
    X"f0", X"90", X"18", X"7b", X"e0", X"a4", X"f8", X"a9", 
    X"f0", X"8a", X"f0", X"e0", X"a4", X"29", X"f9", X"8b", 
    X"f0", X"a3", X"e0", X"a4", X"29", X"f5", X"83", X"88", 
    X"82", X"22", X"22", X"ac", X"82", X"ad", X"83", X"90", 
    X"18", X"7e", X"e0", X"fe", X"a3", X"e0", X"ff", X"be", 
    X"00", X"03", X"60", X"12", X"1f", X"0f", X"90", X"18", 
    X"7d", X"e0", X"8c", X"82", X"8d", X"83", X"12", X"66", 
    X"a0", X"a3", X"de", X"fa", X"df", X"f8", X"8c", X"82", 
    X"8d", X"83", X"22", X"af", X"f0", X"ae", X"83", X"e5", 
    X"82", X"90", X"18", X"85", X"f0", X"ee", X"a3", X"f0", 
    X"ef", X"a3", X"f0", X"90", X"18", X"85", X"e0", X"f5", 
    X"13", X"a3", X"e0", X"f5", X"14", X"a3", X"e0", X"f5", 
    X"15", X"aa", X"13", X"ab", X"14", X"ac", X"15", X"90", 
    X"18", X"80", X"e0", X"f8", X"a3", X"e0", X"f9", X"a3", 
    X"e0", X"ff", X"90", X"18", X"83", X"e0", X"f5", X"16", 
    X"a3", X"e0", X"f5", X"17", X"ad", X"16", X"ae", X"17", 
    X"15", X"16", X"74", X"ff", X"b5", X"16", X"02", X"15", 
    X"17", X"ed", X"4e", X"60", X"20", X"88", X"82", X"89", 
    X"83", X"8f", X"f0", X"12", X"70", X"5a", X"fe", X"a3", 
    X"a8", X"82", X"a9", X"83", X"8a", X"82", X"8b", X"83", 
    X"8c", X"f0", X"ee", X"12", X"66", X"a0", X"a3", X"aa", 
    X"82", X"ab", X"83", X"80", X"cf", X"85", X"13", X"82", 
    X"85", X"14", X"83", X"85", X"15", X"f0", X"22", X"c0", 
    X"0c", X"85", X"81", X"0c", X"7e", X"00", X"8e", X"83", 
    X"12", X"66", X"87", X"d0", X"0c", X"22", X"af", X"f0", 
    X"ae", X"83", X"e5", X"82", X"90", X"18", X"89", X"f0", 
    X"ee", X"a3", X"f0", X"ef", X"a3", X"f0", X"90", X"18", 
    X"89", X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", 
    X"ff", X"90", X"18", X"88", X"e0", X"fc", X"90", X"18", 
    X"9d", X"e4", X"f0", X"a3", X"f0", X"a3", X"f0", X"90", 
    X"18", X"a0", X"ed", X"f0", X"ee", X"a3", X"f0", X"ef", 
    X"a3", X"f0", X"90", X"18", X"a3", X"ec", X"f0", X"90", 
    X"67", X"77", X"02", X"68", X"d5", X"c0", X"0c", X"85", 
    X"81", X"0c", X"e5", X"0c", X"24", X"fb", X"ff", X"90", 
    X"18", X"9d", X"e4", X"f0", X"a3", X"f0", X"a3", X"f0", 
    X"e5", X"0c", X"24", X"fb", X"f8", X"90", X"18", X"a0", 
    X"e6", X"f0", X"08", X"e6", X"a3", X"f0", X"08", X"e6", 
    X"a3", X"f0", X"90", X"18", X"a3", X"ef", X"f0", X"90", 
    X"67", X"77", X"12", X"68", X"d5", X"d0", X"0c", X"22", 
    X"e5", X"82", X"90", X"18", X"99", X"f0", X"e0", X"ff", 
    X"90", X"18", X"8f", X"e0", X"c0", X"e0", X"a3", X"e0", 
    X"c0", X"e0", X"a3", X"e0", X"c0", X"e0", X"12", X"68", 
    X"13", X"80", X"0d", X"90", X"18", X"8d", X"e0", X"c0", 
    X"e0", X"a3", X"e0", X"c0", X"e0", X"8f", X"82", X"22", 
    X"15", X"81", X"15", X"81", X"15", X"81", X"90", X"18", 
    X"97", X"e0", X"24", X"01", X"f0", X"a3", X"e0", X"34", 
    X"00", X"f0", X"22", X"e5", X"82", X"90", X"18", X"9a", 
    X"f0", X"e0", X"24", X"30", X"ff", X"24", X"c6", X"50", 
    X"13", X"74", X"07", X"2f", X"ff", X"90", X"18", X"8c", 
    X"e0", X"60", X"09", X"8f", X"05", X"7e", X"00", X"43", 
    X"05", X"20", X"8d", X"07", X"8f", X"82", X"02", X"67", 
    X"f8", X"e5", X"82", X"90", X"18", X"9b", X"f0", X"e0", 
    X"ff", X"c4", X"54", X"0f", X"f5", X"82", X"c0", X"07", 
    X"12", X"68", X"33", X"d0", X"07", X"53", X"07", X"0f", 
    X"8f", X"82", X"02", X"68", X"33", X"e5", X"82", X"90", 
    X"18", X"9c", X"f0", X"90", X"18", X"92", X"e0", X"fc", 
    X"a3", X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", 
    X"ff", X"90", X"18", X"96", X"e0", X"fb", X"75", X"13", 
    X"20", X"90", X"18", X"9c", X"e0", X"f9", X"8b", X"00", 
    X"e8", X"28", X"f8", X"ef", X"23", X"54", X"01", X"48", 
    X"fb", X"ec", X"2c", X"fc", X"ed", X"33", X"fd", X"ee", 
    X"33", X"fe", X"ef", X"33", X"ff", X"c3", X"eb", X"99", 
    X"40", X"07", X"eb", X"c3", X"99", X"fb", X"43", X"04", 
    X"01", X"e5", X"13", X"14", X"fa", X"8a", X"13", X"70", 
    X"d5", X"90", X"18", X"92", X"ec", X"f0", X"ed", X"a3", 
    X"f0", X"ee", X"a3", X"f0", X"ef", X"a3", X"f0", X"90", 
    X"18", X"96", X"eb", X"f0", X"22", X"af", X"83", X"e5", 
    X"82", X"90", X"18", X"a4", X"f0", X"ef", X"a3", X"f0", 
    X"90", X"18", X"a4", X"e0", X"fe", X"a3", X"e0", X"ff", 
    X"90", X"18", X"8d", X"ee", X"f0", X"ef", X"a3", X"f0", 
    X"90", X"18", X"9d", X"e0", X"fd", X"a3", X"e0", X"fe", 
    X"a3", X"e0", X"ff", X"90", X"18", X"8f", X"ed", X"f0", 
    X"ee", X"a3", X"f0", X"ef", X"a3", X"f0", X"90", X"18", 
    X"97", X"e4", X"f0", X"a3", X"f0", X"90", X"18", X"a0", 
    X"e0", X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", 
    X"8d", X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", 
    X"5a", X"fc", X"90", X"18", X"a0", X"74", X"01", X"2d", 
    X"f0", X"e4", X"3e", X"a3", X"f0", X"ef", X"a3", X"f0", 
    X"ec", X"70", X"03", X"02", X"70", X"36", X"bc", X"25", 
    X"02", X"80", X"03", X"02", X"70", X"2e", X"90", X"18", 
    X"a6", X"e4", X"f0", X"90", X"18", X"a7", X"f0", X"90", 
    X"18", X"a8", X"f0", X"90", X"18", X"a9", X"f0", X"90", 
    X"18", X"aa", X"f0", X"90", X"18", X"ab", X"f0", X"90", 
    X"18", X"ac", X"f0", X"90", X"18", X"ad", X"f0", X"90", 
    X"18", X"af", X"f0", X"90", X"18", X"b0", X"f0", X"90", 
    X"18", X"b1", X"14", X"f0", X"90", X"18", X"a0", X"e0", 
    X"fd", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"8d", 
    X"82", X"8e", X"83", X"8f", X"f0", X"12", X"70", X"5a", 
    X"fb", X"a3", X"ad", X"82", X"ae", X"83", X"90", X"18", 
    X"a0", X"ed", X"f0", X"ee", X"a3", X"f0", X"ef", X"a3", 
    X"f0", X"90", X"18", X"b3", X"eb", X"f0", X"bb", X"25", 
    X"08", X"8b", X"82", X"12", X"67", X"f8", X"02", X"69", 
    X"0d", X"bb", X"30", X"00", X"40", X"43", X"eb", X"24", 
    X"c6", X"40", X"3e", X"90", X"18", X"b1", X"e0", X"fa", 
    X"ba", X"ff", X"27", X"c0", X"05", X"c0", X"06", X"c0", 
    X"07", X"90", X"18", X"b0", X"e0", X"75", X"f0", X"0a", 
    X"a4", X"ff", X"8b", X"06", X"ee", X"2f", X"24", X"d0", 
    X"f0", X"d0", X"07", X"d0", X"06", X"d0", X"05", X"e0", 
    X"70", X"a5", X"90", X"18", X"a7", X"74", X"01", X"f0", 
    X"80", X"9d", X"ea", X"75", X"f0", X"0a", X"a4", X"fa", 
    X"2b", X"24", X"d0", X"90", X"18", X"b1", X"f0", X"80", 
    X"8e", X"90", X"18", X"b3", X"e0", X"fb", X"bb", X"2e", 
    X"15", X"90", X"18", X"b1", X"e0", X"fa", X"ba", X"ff", 
    X"02", X"80", X"03", X"02", X"69", X"77", X"90", X"18", 
    X"b1", X"e4", X"f0", X"02", X"69", X"77", X"bb", X"61", 
    X"00", X"40", X"14", X"eb", X"24", X"85", X"40", X"0f", 
    X"90", X"18", X"b3", X"74", X"df", X"5b", X"f0", X"90", 
    X"18", X"8c", X"74", X"01", X"f0", X"80", X"05", X"90", 
    X"18", X"8c", X"e4", X"f0", X"90", X"18", X"b3", X"e0", 
    X"fb", X"bb", X"20", X"02", X"80", X"75", X"bb", X"2b", 
    X"02", X"80", X"67", X"bb", X"2d", X"02", X"80", X"59", 
    X"bb", X"42", X"02", X"80", X"6f", X"bb", X"43", X"02", 
    X"80", X"7c", X"bb", X"44", X"03", X"02", X"6c", X"7c", 
    X"bb", X"46", X"03", X"02", X"6c", X"a2", X"bb", X"48", 
    X"03", X"02", X"69", X"77", X"bb", X"49", X"03", X"02", 
    X"6c", X"7c", X"bb", X"4a", X"03", X"02", X"69", X"77", 
    X"bb", X"4c", X"02", X"80", X"50", X"bb", X"4f", X"03", 
    X"02", X"6c", X"8a", X"bb", X"50", X"03", X"02", X"6b", 
    X"ed", X"bb", X"53", X"02", X"80", X"77", X"bb", X"54", 
    X"03", X"02", X"69", X"77", X"bb", X"55", X"03", X"02", 
    X"6c", X"92", X"bb", X"58", X"03", X"02", X"6c", X"9a", 
    X"bb", X"5a", X"03", X"02", X"69", X"77", X"02", X"6c", 
    X"aa", X"90", X"18", X"a6", X"74", X"01", X"f0", X"02", 
    X"69", X"77", X"90", X"18", X"a8", X"74", X"01", X"f0", 
    X"02", X"69", X"77", X"90", X"18", X"a9", X"74", X"01", 
    X"f0", X"02", X"69", X"77", X"90", X"18", X"ab", X"74", 
    X"01", X"f0", X"02", X"69", X"77", X"90", X"18", X"ac", 
    X"74", X"01", X"f0", X"02", X"69", X"77", X"90", X"18", 
    X"ab", X"e0", X"60", X"0e", X"90", X"18", X"a3", X"e0", 
    X"14", X"f9", X"f0", X"90", X"18", X"b3", X"e7", X"f0", 
    X"80", X"0f", X"90", X"18", X"a3", X"e0", X"24", X"fe", 
    X"ff", X"f0", X"8f", X"01", X"90", X"18", X"b3", X"e7", 
    X"f0", X"90", X"18", X"b3", X"e0", X"f5", X"82", X"12", 
    X"67", X"f8", X"02", X"6c", X"b6", X"90", X"18", X"a3", 
    X"e0", X"24", X"fd", X"ff", X"f0", X"8f", X"01", X"87", 
    X"05", X"09", X"87", X"06", X"09", X"87", X"07", X"19", 
    X"19", X"90", X"18", X"92", X"ed", X"f0", X"ee", X"a3", 
    X"f0", X"ef", X"a3", X"f0", X"8d", X"82", X"8e", X"83", 
    X"8f", X"f0", X"12", X"70", X"42", X"ae", X"82", X"90", 
    X"18", X"b1", X"e0", X"ff", X"bf", X"ff", X"05", X"90", 
    X"18", X"b1", X"ee", X"f0", X"90", X"18", X"a6", X"e0", 
    X"70", X"2e", X"90", X"18", X"b0", X"e0", X"ff", X"c3", 
    X"ee", X"9f", X"50", X"24", X"90", X"18", X"b0", X"ef", 
    X"c3", X"9e", X"f0", X"e0", X"ff", X"8f", X"05", X"1f", 
    X"ed", X"60", X"10", X"75", X"82", X"20", X"c0", X"07", 
    X"c0", X"06", X"12", X"67", X"f8", X"d0", X"06", X"d0", 
    X"07", X"80", X"ea", X"90", X"18", X"b0", X"ef", X"f0", 
    X"90", X"18", X"b1", X"e0", X"ff", X"c0", X"06", X"90", 
    X"18", X"92", X"e0", X"fa", X"a3", X"e0", X"fd", X"a3", 
    X"e0", X"fe", X"8a", X"82", X"8d", X"83", X"8e", X"f0", 
    X"12", X"70", X"5a", X"f5", X"0d", X"d0", X"06", X"e5", 
    X"0d", X"60", X"3e", X"8f", X"05", X"1f", X"c3", X"74", 
    X"80", X"8d", X"f0", X"63", X"f0", X"80", X"95", X"f0", 
    X"50", X"2f", X"c0", X"06", X"85", X"0d", X"82", X"c0", 
    X"07", X"c0", X"06", X"12", X"67", X"f8", X"d0", X"06", 
    X"d0", X"07", X"90", X"18", X"92", X"e0", X"fa", X"a3", 
    X"e0", X"fd", X"a3", X"e0", X"fe", X"0a", X"ba", X"00", 
    X"01", X"0d", X"90", X"18", X"92", X"ea", X"f0", X"ed", 
    X"a3", X"f0", X"ee", X"a3", X"f0", X"d0", X"06", X"80", 
    X"a4", X"90", X"18", X"a6", X"e0", X"70", X"03", X"02", 
    X"6c", X"b6", X"90", X"18", X"b0", X"e0", X"ff", X"c3", 
    X"ee", X"9f", X"40", X"03", X"02", X"6c", X"b6", X"90", 
    X"18", X"b0", X"ef", X"c3", X"9e", X"f0", X"e0", X"ff", 
    X"8f", X"06", X"1f", X"ee", X"70", X"03", X"02", X"6c", 
    X"b1", X"75", X"82", X"20", X"c0", X"07", X"12", X"67", 
    X"f8", X"d0", X"07", X"80", X"eb", X"90", X"18", X"a3", 
    X"e0", X"24", X"fd", X"fe", X"f0", X"8e", X"01", X"87", 
    X"02", X"09", X"87", X"05", X"09", X"87", X"06", X"19", 
    X"19", X"90", X"18", X"92", X"ea", X"f0", X"ed", X"a3", 
    X"f0", X"ee", X"a3", X"f0", X"90", X"18", X"94", X"e0", 
    X"fe", X"be", X"80", X"00", X"40", X"08", X"90", X"18", 
    X"b3", X"74", X"43", X"f0", X"80", X"20", X"be", X"60", 
    X"00", X"40", X"08", X"90", X"18", X"b3", X"74", X"50", 
    X"f0", X"80", X"13", X"be", X"40", X"00", X"40", X"08", 
    X"90", X"18", X"b3", X"74", X"49", X"f0", X"80", X"06", 
    X"90", X"18", X"b3", X"74", X"58", X"f0", X"90", X"18", 
    X"b3", X"e0", X"fe", X"f5", X"82", X"c0", X"06", X"12", 
    X"67", X"f8", X"75", X"82", X"3a", X"12", X"67", X"f8", 
    X"75", X"82", X"30", X"12", X"67", X"f8", X"75", X"82", 
    X"78", X"12", X"67", X"f8", X"d0", X"06", X"be", X"49", 
    X"02", X"80", X"0e", X"be", X"50", X"02", X"80", X"09", 
    X"90", X"18", X"93", X"e0", X"f5", X"82", X"12", X"68", 
    X"59", X"90", X"18", X"92", X"e0", X"f5", X"82", X"12", 
    X"68", X"59", X"80", X"3a", X"90", X"18", X"aa", X"74", 
    X"01", X"f0", X"90", X"18", X"af", X"74", X"0a", X"f0", 
    X"80", X"2c", X"90", X"18", X"af", X"74", X"08", X"f0", 
    X"80", X"24", X"90", X"18", X"af", X"74", X"0a", X"f0", 
    X"80", X"1c", X"90", X"18", X"af", X"74", X"10", X"f0", 
    X"80", X"14", X"90", X"18", X"ad", X"74", X"01", X"f0", 
    X"80", X"0c", X"8b", X"82", X"12", X"67", X"f8", X"80", 
    X"05", X"90", X"18", X"b0", X"ef", X"f0", X"90", X"18", 
    X"ad", X"e0", X"60", X"71", X"90", X"18", X"a3", X"e0", 
    X"24", X"fc", X"ff", X"f0", X"8f", X"01", X"87", X"03", 
    X"09", X"87", X"05", X"09", X"87", X"06", X"09", X"87", 
    X"07", X"19", X"19", X"19", X"90", X"18", X"92", X"eb", 
    X"f0", X"ed", X"a3", X"f0", X"ee", X"a3", X"f0", X"ef", 
    X"a3", X"f0", X"90", X"18", X"92", X"74", X"f0", X"f0", 
    X"74", X"70", X"a3", X"f0", X"74", X"80", X"a3", X"f0", 
    X"90", X"18", X"92", X"e0", X"f5", X"0e", X"a3", X"e0", 
    X"f5", X"0f", X"a3", X"e0", X"f5", X"10", X"74", X"01", 
    X"25", X"0e", X"fa", X"e4", X"35", X"0f", X"fb", X"af", 
    X"10", X"90", X"18", X"92", X"ea", X"f0", X"eb", X"a3", 
    X"f0", X"ef", X"a3", X"f0", X"85", X"0e", X"82", X"85", 
    X"0f", X"83", X"85", X"10", X"f0", X"12", X"70", X"5a", 
    X"ff", X"70", X"03", X"02", X"69", X"0d", X"8f", X"82", 
    X"12", X"67", X"f8", X"80", X"c3", X"90", X"18", X"af", 
    X"e0", X"70", X"03", X"02", X"69", X"0d", X"90", X"18", 
    X"ab", X"e0", X"60", X"47", X"90", X"18", X"a3", X"e0", 
    X"14", X"f9", X"f0", X"87", X"07", X"7e", X"00", X"7d", 
    X"00", X"7b", X"00", X"90", X"18", X"92", X"ef", X"f0", 
    X"ee", X"a3", X"f0", X"ed", X"a3", X"f0", X"eb", X"a3", 
    X"f0", X"90", X"18", X"aa", X"e0", X"60", X"03", X"02", 
    X"6d", X"f9", X"90", X"18", X"92", X"e0", X"fb", X"a3", 
    X"e0", X"a3", X"e0", X"a3", X"e0", X"7d", X"00", X"7e", 
    X"00", X"7f", X"00", X"90", X"18", X"92", X"eb", X"f0", 
    X"ed", X"a3", X"f0", X"ee", X"a3", X"f0", X"ef", X"a3", 
    X"f0", X"80", X"76", X"90", X"18", X"ac", X"e0", X"60", 
    X"28", X"90", X"18", X"a3", X"e0", X"24", X"fc", X"ff", 
    X"f0", X"8f", X"01", X"87", X"03", X"09", X"87", X"05", 
    X"09", X"87", X"06", X"09", X"87", X"07", X"19", X"19", 
    X"19", X"90", X"18", X"92", X"eb", X"f0", X"ed", X"a3", 
    X"f0", X"ee", X"a3", X"f0", X"ef", X"a3", X"f0", X"80", 
    X"48", X"90", X"18", X"a3", X"e0", X"24", X"fe", X"ff", 
    X"f0", X"8f", X"01", X"87", X"06", X"09", X"87", X"07", 
    X"19", X"ef", X"33", X"95", X"e0", X"fd", X"fb", X"90", 
    X"18", X"92", X"ee", X"f0", X"ef", X"a3", X"f0", X"ed", 
    X"a3", X"f0", X"eb", X"a3", X"f0", X"90", X"18", X"aa", 
    X"e0", X"70", X"1e", X"90", X"18", X"92", X"e0", X"fb", 
    X"a3", X"e0", X"fd", X"a3", X"e0", X"a3", X"e0", X"7e", 
    X"00", X"7f", X"00", X"90", X"18", X"92", X"eb", X"f0", 
    X"ed", X"a3", X"f0", X"ee", X"a3", X"f0", X"ef", X"a3", 
    X"f0", X"90", X"18", X"aa", X"e0", X"60", X"41", X"90", 
    X"18", X"92", X"e0", X"fb", X"a3", X"e0", X"fd", X"a3", 
    X"e0", X"fe", X"a3", X"e0", X"ff", X"30", X"e7", X"2b", 
    X"90", X"18", X"92", X"e0", X"fb", X"a3", X"e0", X"fd", 
    X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"c3", X"e4", 
    X"9b", X"fb", X"e4", X"9d", X"fd", X"e4", X"9e", X"fe", 
    X"e4", X"9f", X"ff", X"90", X"18", X"92", X"eb", X"f0", 
    X"ed", X"a3", X"f0", X"ee", X"a3", X"f0", X"ef", X"a3", 
    X"f0", X"80", X"05", X"90", X"18", X"aa", X"e4", X"f0", 
    X"90", X"18", X"ae", X"74", X"01", X"f0", X"90", X"18", 
    X"af", X"e0", X"f5", X"0e", X"75", X"11", X"b9", X"75", 
    X"12", X"18", X"75", X"0d", X"00", X"90", X"18", X"96", 
    X"e4", X"f0", X"85", X"0e", X"82", X"12", X"68", X"75", 
    X"90", X"18", X"ae", X"e0", X"70", X"23", X"90", X"18", 
    X"96", X"e0", X"c4", X"fa", X"85", X"11", X"82", X"85", 
    X"12", X"83", X"e0", X"ff", X"42", X"02", X"85", X"11", 
    X"82", X"85", X"12", X"83", X"ea", X"f0", X"15", X"11", 
    X"74", X"ff", X"b5", X"11", X"02", X"15", X"12", X"80", 
    X"0c", X"90", X"18", X"96", X"e0", X"fa", X"85", X"11", 
    X"82", X"85", X"12", X"83", X"f0", X"05", X"0d", X"90", 
    X"18", X"ae", X"e0", X"b4", X"01", X"00", X"e4", X"33", 
    X"f0", X"90", X"18", X"92", X"e0", X"fa", X"a3", X"e0", 
    X"fb", X"a3", X"e0", X"fe", X"a3", X"e0", X"ff", X"ea", 
    X"4b", X"4e", X"4f", X"70", X"a0", X"90", X"18", X"ba", 
    X"e5", X"11", X"f0", X"e5", X"12", X"a3", X"f0", X"90", 
    X"18", X"b2", X"e5", X"0d", X"f0", X"90", X"18", X"b0", 
    X"e0", X"70", X"06", X"90", X"18", X"b0", X"74", X"01", 
    X"f0", X"90", X"18", X"a7", X"e0", X"ff", X"e0", X"70", 
    X"2f", X"90", X"18", X"a6", X"e0", X"70", X"29", X"ae", 
    X"0d", X"90", X"18", X"b0", X"e0", X"fd", X"8e", X"03", 
    X"0b", X"c3", X"eb", X"9d", X"50", X"15", X"75", X"82", 
    X"20", X"c0", X"07", X"c0", X"06", X"c0", X"05", X"12", 
    X"67", X"f8", X"d0", X"05", X"d0", X"06", X"d0", X"07", 
    X"1d", X"80", X"e3", X"90", X"18", X"b0", X"ed", X"f0", 
    X"90", X"18", X"aa", X"e0", X"60", X"12", X"75", X"82", 
    X"2d", X"c0", X"07", X"12", X"67", X"f8", X"d0", X"07", 
    X"90", X"18", X"b0", X"e0", X"14", X"f0", X"80", X"34", 
    X"90", X"18", X"b2", X"e0", X"60", X"2e", X"90", X"18", 
    X"a8", X"e0", X"60", X"12", X"75", X"82", X"2b", X"c0", 
    X"07", X"12", X"67", X"f8", X"d0", X"07", X"90", X"18", 
    X"b0", X"e0", X"14", X"f0", X"80", X"16", X"90", X"18", 
    X"a9", X"e0", X"60", X"10", X"75", X"82", X"20", X"c0", 
    X"07", X"12", X"67", X"f8", X"d0", X"07", X"90", X"18", 
    X"b0", X"e0", X"14", X"f0", X"90", X"18", X"a6", X"e0", 
    X"70", X"32", X"90", X"18", X"b2", X"e0", X"fe", X"90", 
    X"18", X"b0", X"e0", X"fd", X"8d", X"03", X"1d", X"c3", 
    X"ee", X"9b", X"50", X"3e", X"ef", X"60", X"06", X"7a", 
    X"30", X"7b", X"00", X"80", X"04", X"7a", X"20", X"7b", 
    X"00", X"8a", X"82", X"c0", X"07", X"c0", X"06", X"c0", 
    X"05", X"12", X"67", X"f8", X"d0", X"05", X"d0", X"06", 
    X"d0", X"07", X"80", X"d8", X"90", X"18", X"b0", X"e0", 
    X"ff", X"90", X"18", X"b2", X"e0", X"fe", X"c3", X"9f", 
    X"50", X"09", X"90", X"18", X"b0", X"ef", X"c3", X"9e", 
    X"f0", X"80", X"0c", X"90", X"18", X"b0", X"e4", X"f0", 
    X"80", X"05", X"90", X"18", X"b0", X"ed", X"f0", X"90", 
    X"18", X"ba", X"e0", X"fe", X"a3", X"e0", X"ff", X"90", 
    X"18", X"b2", X"e0", X"fd", X"8d", X"03", X"1d", X"eb", 
    X"60", X"49", X"90", X"18", X"ae", X"e0", X"b4", X"01", 
    X"00", X"e4", X"33", X"f0", X"90", X"18", X"ae", X"e0", 
    X"70", X"14", X"0e", X"be", X"00", X"01", X"0f", X"8e", 
    X"82", X"8f", X"83", X"e0", X"c4", X"54", X"0f", X"fb", 
    X"90", X"18", X"96", X"f0", X"80", X"0e", X"8e", X"82", 
    X"8f", X"83", X"e0", X"fb", X"53", X"03", X"0f", X"90", 
    X"18", X"96", X"eb", X"f0", X"90", X"18", X"96", X"e0", 
    X"f5", X"82", X"c0", X"07", X"c0", X"06", X"c0", X"05", 
    X"12", X"68", X"33", X"d0", X"05", X"d0", X"06", X"d0", 
    X"07", X"80", X"b1", X"90", X"18", X"a6", X"e0", X"70", 
    X"03", X"02", X"69", X"0d", X"90", X"18", X"b0", X"e0", 
    X"ff", X"8f", X"06", X"1f", X"ee", X"70", X"03", X"02", 
    X"69", X"0d", X"75", X"82", X"20", X"c0", X"07", X"12", 
    X"67", X"f8", X"d0", X"07", X"80", X"eb", X"8c", X"82", 
    X"12", X"67", X"f8", X"02", X"69", X"0d", X"90", X"18", 
    X"97", X"e0", X"fe", X"a3", X"e0", X"8e", X"82", X"f5", 
    X"83", X"22", X"aa", X"82", X"ab", X"83", X"12", X"70", 
    X"5a", X"60", X"03", X"a3", X"80", X"f8", X"c3", X"e5", 
    X"82", X"9a", X"f5", X"82", X"e5", X"83", X"9b", X"f5", 
    X"83", X"22", X"20", X"f7", X"14", X"30", X"f6", X"14", 
    X"88", X"83", X"a8", X"82", X"20", X"f5", X"07", X"e6", 
    X"a8", X"83", X"75", X"83", X"00", X"22", X"e2", X"80", 
    X"f7", X"e4", X"93", X"22", X"e0", X"22", X"75", X"82", 
    X"00", X"22", X"54", X"61", X"73", X"6b", X"20", X"31", 
    X"00", X"54", X"61", X"73", X"6b", X"20", X"32", X"00", 
    X"0a", X"0d", X"00", X"4c", X"69", X"67", X"68", X"74", 
    X"35", X"32", X"20", X"70", X"72", X"6f", X"6a", X"65", 
    X"63", X"74", X"20", X"2d", X"2d", X"20", X"4e", X"6f", 
    X"76", X"20", X"20", X"32", X"20", X"32", X"30", X"31", 
    X"38", X"20", X"31", X"37", X"3a", X"31", X"38", X"3a", 
    X"31", X"37", X"0a", X"0a", X"0d", X"00", X"46", X"72", 
    X"65", X"65", X"52", X"54", X"4f", X"53", X"20", X"74", 
    X"65", X"73", X"74", X"2e", X"0a", X"0d", X"00", X"42", 
    X"6c", X"69", X"6e", X"6b", X"54", X"61", X"73", X"6b", 
    X"00", X"52", X"58", X"54", X"61", X"73", X"6b", X"00", 
    X"48", X"61", X"6c", X"6c", X"6f", X"20", X"76", X"6f", 
    X"6e", X"20", X"25", X"73", X"21", X"0a", X"0d", X"00", 
    X"25", X"63", X"00", X"49", X"44", X"4c", X"45", X"00", 
    X"3c", X"4e", X"4f", X"20", X"46", X"4c", X"4f", X"41", 
    X"54", X"3e", X"00" 
);


end package obj_code_pkg;
